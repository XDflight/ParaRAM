magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -465 23 465 42
rect -465 -23 -446 23
rect 446 -23 465 23
rect -465 -42 465 -23
<< polycontact >>
rect -446 -23 446 23
<< metal1 >>
rect -457 23 457 34
rect -457 -23 -446 23
rect 446 -23 457 23
rect -457 -34 457 -23
<< properties >>
string GDS_END 659484
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 658712
<< end >>
