magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 348
<< mvpmos >>
rect 0 0 120 228
rect 224 0 344 228
<< mvpdiff >>
rect -88 215 0 228
rect -88 169 -75 215
rect -29 169 0 215
rect -88 59 0 169
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 215 224 228
rect 120 169 149 215
rect 195 169 224 215
rect 120 59 224 169
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 215 432 228
rect 344 169 373 215
rect 419 169 432 215
rect 344 59 432 169
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 169 -29 215
rect -75 13 -29 59
rect 149 169 195 215
rect 149 13 195 59
rect 373 169 419 215
rect 373 13 419 59
<< polysilicon >>
rect 0 228 120 272
rect 224 228 344 272
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 215 -29 228
rect -75 59 -29 169
rect -75 0 -29 13
rect 149 215 195 228
rect 149 59 195 169
rect 149 0 195 13
rect 373 215 419 228
rect 373 59 419 169
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 114 -52 114 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 114 396 114 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 114 172 114 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 118000
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 116274
<< end >>
