magic
tech gf180mcuB
timestamp 1667403374
<< metal1 >>
rect 0 147 44 159
rect 11 106 16 147
rect 28 99 33 140
rect 26 93 36 99
rect 28 92 33 93
rect 11 9 16 33
rect 0 -3 44 9
<< obsm1 >>
rect 23 41 33 46
rect 28 16 33 41
<< metal2 >>
rect 10 154 18 155
rect 9 148 19 154
rect 10 147 18 148
rect 26 92 36 100
rect 10 8 18 9
rect 9 2 19 8
rect 10 1 18 2
<< labels >>
rlabel metal2 s 10 147 18 155 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 147 44 159 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 2 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 2 nsew ground bidirectional
rlabel metal1 s 0 -3 44 9 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 26 92 36 100 6 Y
port 3 nsew signal output
rlabel metal1 s 28 92 33 140 6 Y
port 3 nsew signal output
rlabel metal1 s 26 93 36 99 6 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 44 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
