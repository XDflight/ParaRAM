magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 7030 1094
<< pwell >>
rect -86 -86 7030 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 1916 69 2036 333
rect 2140 69 2260 333
rect 2364 69 2484 333
rect 2588 69 2708 333
rect 2812 69 2932 333
rect 3036 69 3156 333
rect 3260 69 3380 333
rect 3484 69 3604 333
rect 3708 69 3828 333
rect 3932 69 4052 333
rect 4156 69 4276 333
rect 4380 69 4500 333
rect 4604 69 4724 333
rect 4828 69 4948 333
rect 5052 69 5172 333
rect 5276 69 5396 333
rect 5500 69 5620 333
rect 5724 69 5844 333
rect 5948 69 6068 333
rect 6172 69 6292 333
rect 6396 69 6516 333
rect 6620 69 6740 333
<< mvpmos >>
rect 124 573 224 939
rect 348 573 448 939
rect 572 573 672 939
rect 796 573 896 939
rect 1020 573 1120 939
rect 1244 573 1344 939
rect 1468 573 1568 939
rect 1692 573 1792 939
rect 1916 573 2016 939
rect 2140 573 2240 939
rect 2364 573 2464 939
rect 2588 573 2688 939
rect 2812 573 2912 939
rect 3036 573 3136 939
rect 3260 573 3360 939
rect 3484 573 3584 939
rect 3708 573 3808 939
rect 3932 573 4032 939
rect 4156 573 4256 939
rect 4380 573 4480 939
rect 4604 573 4704 939
rect 4828 573 4928 939
rect 5052 573 5152 939
rect 5276 573 5376 939
rect 5500 573 5600 939
rect 5724 573 5824 939
rect 5948 573 6048 939
rect 6172 573 6272 939
rect 6396 573 6496 939
rect 6620 573 6720 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 244 287 348 333
rect 244 147 273 287
rect 319 147 348 287
rect 244 69 348 147
rect 468 287 572 333
rect 468 147 497 287
rect 543 147 572 287
rect 468 69 572 147
rect 692 287 796 333
rect 692 147 721 287
rect 767 147 796 287
rect 692 69 796 147
rect 916 287 1020 333
rect 916 147 945 287
rect 991 147 1020 287
rect 916 69 1020 147
rect 1140 287 1244 333
rect 1140 147 1169 287
rect 1215 147 1244 287
rect 1140 69 1244 147
rect 1364 287 1468 333
rect 1364 147 1393 287
rect 1439 147 1468 287
rect 1364 69 1468 147
rect 1588 287 1692 333
rect 1588 147 1617 287
rect 1663 147 1692 287
rect 1588 69 1692 147
rect 1812 287 1916 333
rect 1812 147 1841 287
rect 1887 147 1916 287
rect 1812 69 1916 147
rect 2036 287 2140 333
rect 2036 147 2065 287
rect 2111 147 2140 287
rect 2036 69 2140 147
rect 2260 287 2364 333
rect 2260 147 2289 287
rect 2335 147 2364 287
rect 2260 69 2364 147
rect 2484 287 2588 333
rect 2484 147 2513 287
rect 2559 147 2588 287
rect 2484 69 2588 147
rect 2708 287 2812 333
rect 2708 147 2737 287
rect 2783 147 2812 287
rect 2708 69 2812 147
rect 2932 287 3036 333
rect 2932 147 2961 287
rect 3007 147 3036 287
rect 2932 69 3036 147
rect 3156 287 3260 333
rect 3156 147 3185 287
rect 3231 147 3260 287
rect 3156 69 3260 147
rect 3380 287 3484 333
rect 3380 147 3409 287
rect 3455 147 3484 287
rect 3380 69 3484 147
rect 3604 287 3708 333
rect 3604 147 3633 287
rect 3679 147 3708 287
rect 3604 69 3708 147
rect 3828 287 3932 333
rect 3828 147 3857 287
rect 3903 147 3932 287
rect 3828 69 3932 147
rect 4052 287 4156 333
rect 4052 147 4081 287
rect 4127 147 4156 287
rect 4052 69 4156 147
rect 4276 287 4380 333
rect 4276 147 4305 287
rect 4351 147 4380 287
rect 4276 69 4380 147
rect 4500 287 4604 333
rect 4500 147 4529 287
rect 4575 147 4604 287
rect 4500 69 4604 147
rect 4724 287 4828 333
rect 4724 147 4753 287
rect 4799 147 4828 287
rect 4724 69 4828 147
rect 4948 287 5052 333
rect 4948 147 4977 287
rect 5023 147 5052 287
rect 4948 69 5052 147
rect 5172 287 5276 333
rect 5172 147 5201 287
rect 5247 147 5276 287
rect 5172 69 5276 147
rect 5396 287 5500 333
rect 5396 147 5425 287
rect 5471 147 5500 287
rect 5396 69 5500 147
rect 5620 287 5724 333
rect 5620 147 5649 287
rect 5695 147 5724 287
rect 5620 69 5724 147
rect 5844 287 5948 333
rect 5844 147 5873 287
rect 5919 147 5948 287
rect 5844 69 5948 147
rect 6068 287 6172 333
rect 6068 147 6097 287
rect 6143 147 6172 287
rect 6068 69 6172 147
rect 6292 287 6396 333
rect 6292 147 6321 287
rect 6367 147 6396 287
rect 6292 69 6396 147
rect 6516 287 6620 333
rect 6516 147 6545 287
rect 6591 147 6620 287
rect 6516 69 6620 147
rect 6740 287 6828 333
rect 6740 147 6769 287
rect 6815 147 6828 287
rect 6740 69 6828 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 224 861 348 939
rect 224 721 273 861
rect 319 721 348 861
rect 224 573 348 721
rect 448 861 572 939
rect 448 721 477 861
rect 523 721 572 861
rect 448 573 572 721
rect 672 861 796 939
rect 672 721 701 861
rect 747 721 796 861
rect 672 573 796 721
rect 896 861 1020 939
rect 896 721 925 861
rect 971 721 1020 861
rect 896 573 1020 721
rect 1120 861 1244 939
rect 1120 721 1149 861
rect 1195 721 1244 861
rect 1120 573 1244 721
rect 1344 861 1468 939
rect 1344 721 1373 861
rect 1419 721 1468 861
rect 1344 573 1468 721
rect 1568 861 1692 939
rect 1568 721 1597 861
rect 1643 721 1692 861
rect 1568 573 1692 721
rect 1792 861 1916 939
rect 1792 721 1821 861
rect 1867 721 1916 861
rect 1792 573 1916 721
rect 2016 861 2140 939
rect 2016 721 2045 861
rect 2091 721 2140 861
rect 2016 573 2140 721
rect 2240 926 2364 939
rect 2240 786 2269 926
rect 2315 786 2364 926
rect 2240 573 2364 786
rect 2464 861 2588 939
rect 2464 721 2513 861
rect 2559 721 2588 861
rect 2464 573 2588 721
rect 2688 861 2812 939
rect 2688 721 2717 861
rect 2763 721 2812 861
rect 2688 573 2812 721
rect 2912 861 3036 939
rect 2912 721 2941 861
rect 2987 721 3036 861
rect 2912 573 3036 721
rect 3136 861 3260 939
rect 3136 721 3165 861
rect 3211 721 3260 861
rect 3136 573 3260 721
rect 3360 861 3484 939
rect 3360 721 3389 861
rect 3435 721 3484 861
rect 3360 573 3484 721
rect 3584 861 3708 939
rect 3584 721 3613 861
rect 3659 721 3708 861
rect 3584 573 3708 721
rect 3808 861 3932 939
rect 3808 721 3837 861
rect 3883 721 3932 861
rect 3808 573 3932 721
rect 4032 861 4156 939
rect 4032 721 4061 861
rect 4107 721 4156 861
rect 4032 573 4156 721
rect 4256 861 4380 939
rect 4256 721 4285 861
rect 4331 721 4380 861
rect 4256 573 4380 721
rect 4480 861 4604 939
rect 4480 721 4509 861
rect 4555 721 4604 861
rect 4480 573 4604 721
rect 4704 861 4828 939
rect 4704 721 4733 861
rect 4779 721 4828 861
rect 4704 573 4828 721
rect 4928 861 5052 939
rect 4928 721 4957 861
rect 5003 721 5052 861
rect 4928 573 5052 721
rect 5152 861 5276 939
rect 5152 721 5181 861
rect 5227 721 5276 861
rect 5152 573 5276 721
rect 5376 861 5500 939
rect 5376 721 5405 861
rect 5451 721 5500 861
rect 5376 573 5500 721
rect 5600 861 5724 939
rect 5600 721 5629 861
rect 5675 721 5724 861
rect 5600 573 5724 721
rect 5824 861 5948 939
rect 5824 721 5853 861
rect 5899 721 5948 861
rect 5824 573 5948 721
rect 6048 861 6172 939
rect 6048 721 6077 861
rect 6123 721 6172 861
rect 6048 573 6172 721
rect 6272 861 6396 939
rect 6272 721 6301 861
rect 6347 721 6396 861
rect 6272 573 6396 721
rect 6496 861 6620 939
rect 6496 721 6525 861
rect 6571 721 6620 861
rect 6496 573 6620 721
rect 6720 861 6808 939
rect 6720 721 6749 861
rect 6795 721 6808 861
rect 6720 573 6808 721
<< mvndiffc >>
rect 49 147 95 287
rect 273 147 319 287
rect 497 147 543 287
rect 721 147 767 287
rect 945 147 991 287
rect 1169 147 1215 287
rect 1393 147 1439 287
rect 1617 147 1663 287
rect 1841 147 1887 287
rect 2065 147 2111 287
rect 2289 147 2335 287
rect 2513 147 2559 287
rect 2737 147 2783 287
rect 2961 147 3007 287
rect 3185 147 3231 287
rect 3409 147 3455 287
rect 3633 147 3679 287
rect 3857 147 3903 287
rect 4081 147 4127 287
rect 4305 147 4351 287
rect 4529 147 4575 287
rect 4753 147 4799 287
rect 4977 147 5023 287
rect 5201 147 5247 287
rect 5425 147 5471 287
rect 5649 147 5695 287
rect 5873 147 5919 287
rect 6097 147 6143 287
rect 6321 147 6367 287
rect 6545 147 6591 287
rect 6769 147 6815 287
<< mvpdiffc >>
rect 49 721 95 861
rect 273 721 319 861
rect 477 721 523 861
rect 701 721 747 861
rect 925 721 971 861
rect 1149 721 1195 861
rect 1373 721 1419 861
rect 1597 721 1643 861
rect 1821 721 1867 861
rect 2045 721 2091 861
rect 2269 786 2315 926
rect 2513 721 2559 861
rect 2717 721 2763 861
rect 2941 721 2987 861
rect 3165 721 3211 861
rect 3389 721 3435 861
rect 3613 721 3659 861
rect 3837 721 3883 861
rect 4061 721 4107 861
rect 4285 721 4331 861
rect 4509 721 4555 861
rect 4733 721 4779 861
rect 4957 721 5003 861
rect 5181 721 5227 861
rect 5405 721 5451 861
rect 5629 721 5675 861
rect 5853 721 5899 861
rect 6077 721 6123 861
rect 6301 721 6347 861
rect 6525 721 6571 861
rect 6749 721 6795 861
<< polysilicon >>
rect 124 939 224 983
rect 348 939 448 983
rect 572 939 672 983
rect 796 939 896 983
rect 1020 939 1120 983
rect 1244 939 1344 983
rect 1468 939 1568 983
rect 1692 939 1792 983
rect 1916 939 2016 983
rect 2140 939 2240 983
rect 2364 939 2464 983
rect 2588 939 2688 983
rect 2812 939 2912 983
rect 3036 939 3136 983
rect 3260 939 3360 983
rect 3484 939 3584 983
rect 3708 939 3808 983
rect 3932 939 4032 983
rect 4156 939 4256 983
rect 4380 939 4480 983
rect 4604 939 4704 983
rect 4828 939 4928 983
rect 5052 939 5152 983
rect 5276 939 5376 983
rect 5500 939 5600 983
rect 5724 939 5824 983
rect 5948 939 6048 983
rect 6172 939 6272 983
rect 6396 939 6496 983
rect 6620 939 6720 983
rect 124 513 224 573
rect 348 513 448 573
rect 572 513 672 573
rect 796 513 896 573
rect 1020 513 1120 573
rect 1244 513 1344 573
rect 1468 513 1568 573
rect 1692 513 1792 573
rect 1916 513 2016 573
rect 2140 513 2240 573
rect 124 500 2240 513
rect 124 454 137 500
rect 1969 454 2240 500
rect 124 443 2240 454
rect 124 441 2036 443
rect 124 333 244 441
rect 348 333 468 441
rect 572 333 692 441
rect 796 333 916 441
rect 1020 333 1140 441
rect 1244 333 1364 441
rect 1468 333 1588 441
rect 1692 333 1812 441
rect 1916 333 2036 441
rect 2140 377 2240 443
rect 2364 513 2464 573
rect 2588 513 2688 573
rect 2812 513 2912 573
rect 3036 513 3136 573
rect 3260 513 3360 573
rect 3484 513 3584 573
rect 3708 513 3808 573
rect 3932 513 4032 573
rect 4156 513 4256 573
rect 2364 510 4256 513
rect 4380 513 4480 573
rect 4604 513 4704 573
rect 4828 513 4928 573
rect 5052 513 5152 573
rect 5276 513 5376 573
rect 5500 513 5600 573
rect 5724 513 5824 573
rect 5948 513 6048 573
rect 6172 513 6272 573
rect 6396 513 6496 573
rect 4380 510 6496 513
rect 2364 507 6496 510
rect 6620 507 6720 573
rect 2364 500 6720 507
rect 2364 454 2377 500
rect 4209 454 4653 500
rect 6485 454 6720 500
rect 2364 441 6720 454
rect 2140 333 2260 377
rect 2364 333 2484 441
rect 2588 333 2708 441
rect 2812 333 2932 441
rect 3036 333 3156 441
rect 3260 333 3380 441
rect 3484 333 3604 441
rect 3708 333 3828 441
rect 3932 333 4052 441
rect 4156 439 4724 441
rect 4156 333 4276 439
rect 4380 435 4724 439
rect 4380 333 4500 435
rect 4604 333 4724 435
rect 4828 333 4948 441
rect 5052 333 5172 441
rect 5276 333 5396 441
rect 5500 333 5620 441
rect 5724 333 5844 441
rect 5948 333 6068 441
rect 6172 333 6292 441
rect 6396 440 6720 441
rect 6396 333 6516 440
rect 6620 377 6720 440
rect 6620 333 6740 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 1916 25 2036 69
rect 2140 25 2260 69
rect 2364 25 2484 69
rect 2588 25 2708 69
rect 2812 25 2932 69
rect 3036 25 3156 69
rect 3260 25 3380 69
rect 3484 25 3604 69
rect 3708 25 3828 69
rect 3932 25 4052 69
rect 4156 25 4276 69
rect 4380 25 4500 69
rect 4604 25 4724 69
rect 4828 25 4948 69
rect 5052 25 5172 69
rect 5276 25 5396 69
rect 5500 25 5620 69
rect 5724 25 5844 69
rect 5948 25 6068 69
rect 6172 25 6292 69
rect 6396 25 6516 69
rect 6620 25 6740 69
<< polycontact >>
rect 137 454 1969 500
rect 2377 454 4209 500
rect 4653 454 6485 500
<< metal1 >>
rect 0 926 6944 1098
rect 0 918 2269 926
rect 49 861 95 918
rect 49 710 95 721
rect 273 861 319 872
rect 273 664 319 721
rect 477 861 523 918
rect 477 710 523 721
rect 701 861 747 872
rect 701 664 747 721
rect 925 861 971 918
rect 925 710 971 721
rect 1149 861 1195 872
rect 1149 664 1195 721
rect 1373 861 1419 918
rect 1373 710 1419 721
rect 1597 861 1643 872
rect 1597 664 1643 721
rect 1821 861 1867 918
rect 1821 710 1867 721
rect 2045 861 2111 872
rect 2091 721 2111 861
rect 2315 918 6944 926
rect 2269 775 2315 786
rect 2513 861 2559 872
rect 2045 664 2111 721
rect 273 580 2111 664
rect 2045 530 2111 580
rect 2513 664 2559 721
rect 2717 861 2763 918
rect 2717 710 2763 721
rect 2941 861 2987 872
rect 2941 664 2987 721
rect 3165 861 3211 918
rect 3165 710 3211 721
rect 3389 861 3435 872
rect 3389 664 3435 721
rect 3613 861 3659 918
rect 3613 710 3659 721
rect 3837 861 3883 872
rect 3837 664 3883 721
rect 4061 861 4107 918
rect 4061 710 4107 721
rect 4285 861 4331 872
rect 4285 664 4331 721
rect 4509 861 4555 918
rect 4509 710 4555 721
rect 4733 861 4779 872
rect 4733 664 4779 721
rect 4957 861 5003 918
rect 4957 710 5003 721
rect 5181 861 5227 872
rect 5181 664 5227 721
rect 5405 861 5451 918
rect 5405 710 5451 721
rect 5629 861 5675 872
rect 5629 664 5675 721
rect 5853 861 5899 918
rect 5853 710 5899 721
rect 6077 861 6123 872
rect 6077 664 6123 721
rect 6301 861 6347 918
rect 6301 710 6347 721
rect 6525 861 6571 872
rect 6525 664 6571 721
rect 6749 861 6795 918
rect 6749 710 6795 721
rect 2513 577 6571 664
rect 4457 576 6571 577
rect 137 500 1969 530
rect 137 443 1969 454
rect 2045 500 4220 530
rect 2045 454 2377 500
rect 4209 454 4220 500
rect 2045 395 2111 454
rect 4457 406 4607 576
rect 4653 500 6485 530
rect 4653 443 6485 454
rect 273 344 2111 395
rect 49 287 95 298
rect 49 90 95 147
rect 273 287 319 344
rect 273 136 319 147
rect 497 287 543 298
rect 497 90 543 147
rect 721 287 767 344
rect 721 136 767 147
rect 945 287 991 298
rect 945 90 991 147
rect 1169 287 1215 344
rect 1169 136 1215 147
rect 1393 287 1439 298
rect 1393 90 1439 147
rect 1617 287 1663 344
rect 1617 136 1663 147
rect 1841 287 1887 298
rect 1841 90 1887 147
rect 2065 287 2111 344
rect 2513 396 4607 406
rect 2513 344 6591 396
rect 2065 136 2111 147
rect 2289 287 2335 298
rect 2289 90 2335 147
rect 2513 287 2565 344
rect 2559 147 2565 287
rect 2513 136 2565 147
rect 2737 287 2783 298
rect 2737 90 2783 147
rect 2961 287 3007 344
rect 2961 136 3007 147
rect 3185 287 3231 298
rect 3185 90 3231 147
rect 3409 287 3455 344
rect 3409 136 3455 147
rect 3633 287 3679 298
rect 3633 90 3679 147
rect 3857 287 3903 344
rect 3857 136 3903 147
rect 4081 287 4127 298
rect 4081 90 4127 147
rect 4305 287 4351 344
rect 4305 136 4351 147
rect 4529 287 4575 298
rect 4529 90 4575 147
rect 4753 287 4799 344
rect 4753 136 4799 147
rect 4977 287 5023 298
rect 4977 90 5023 147
rect 5201 287 5247 344
rect 5201 136 5247 147
rect 5425 287 5471 298
rect 5425 90 5471 147
rect 5649 287 5695 344
rect 5649 136 5695 147
rect 5873 287 5919 298
rect 5873 90 5919 147
rect 6097 287 6143 344
rect 6097 136 6143 147
rect 6321 287 6367 298
rect 6321 90 6367 147
rect 6545 287 6591 344
rect 6545 136 6591 147
rect 6769 287 6815 298
rect 6769 90 6815 147
rect 0 -90 6944 90
<< labels >>
flabel metal1 s 137 443 1969 530 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 6944 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 6769 90 6815 298 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 6525 664 6571 872 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 6077 664 6123 872 1 Z
port 2 nsew default output
rlabel metal1 s 5629 664 5675 872 1 Z
port 2 nsew default output
rlabel metal1 s 5181 664 5227 872 1 Z
port 2 nsew default output
rlabel metal1 s 4733 664 4779 872 1 Z
port 2 nsew default output
rlabel metal1 s 4285 664 4331 872 1 Z
port 2 nsew default output
rlabel metal1 s 3837 664 3883 872 1 Z
port 2 nsew default output
rlabel metal1 s 3389 664 3435 872 1 Z
port 2 nsew default output
rlabel metal1 s 2941 664 2987 872 1 Z
port 2 nsew default output
rlabel metal1 s 2513 664 2559 872 1 Z
port 2 nsew default output
rlabel metal1 s 2513 577 6571 664 1 Z
port 2 nsew default output
rlabel metal1 s 4457 576 6571 577 1 Z
port 2 nsew default output
rlabel metal1 s 4457 406 4607 576 1 Z
port 2 nsew default output
rlabel metal1 s 2513 396 4607 406 1 Z
port 2 nsew default output
rlabel metal1 s 2513 344 6591 396 1 Z
port 2 nsew default output
rlabel metal1 s 6545 136 6591 344 1 Z
port 2 nsew default output
rlabel metal1 s 6097 136 6143 344 1 Z
port 2 nsew default output
rlabel metal1 s 5649 136 5695 344 1 Z
port 2 nsew default output
rlabel metal1 s 5201 136 5247 344 1 Z
port 2 nsew default output
rlabel metal1 s 4753 136 4799 344 1 Z
port 2 nsew default output
rlabel metal1 s 4305 136 4351 344 1 Z
port 2 nsew default output
rlabel metal1 s 3857 136 3903 344 1 Z
port 2 nsew default output
rlabel metal1 s 3409 136 3455 344 1 Z
port 2 nsew default output
rlabel metal1 s 2961 136 3007 344 1 Z
port 2 nsew default output
rlabel metal1 s 2513 136 2565 344 1 Z
port 2 nsew default output
rlabel metal1 s 6749 775 6795 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6301 775 6347 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5853 775 5899 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 775 5451 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 775 5003 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 775 4555 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 775 4107 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 775 3659 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 775 3211 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 775 2763 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 775 2315 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 775 1867 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 775 1419 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 775 971 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 775 523 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 775 95 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6749 710 6795 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6301 710 6347 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5853 710 5899 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 710 5451 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 710 5003 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 710 4555 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 710 4107 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 710 3659 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 710 3211 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 710 2763 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 710 1867 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 710 1419 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 710 971 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 710 523 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 710 95 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 6321 90 6367 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5873 90 5919 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5425 90 5471 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4977 90 5023 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4529 90 4575 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4081 90 4127 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3633 90 3679 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3185 90 3231 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2737 90 2783 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2289 90 2335 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1841 90 1887 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1393 90 1439 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 6944 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6944 1008
string GDS_END 1299994
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1282740
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
