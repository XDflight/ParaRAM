magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 522
rect 224 0 344 522
<< mvndiff >>
rect -88 509 0 522
rect -88 463 -75 509
rect -29 463 0 509
rect -88 397 0 463
rect -88 351 -75 397
rect -29 351 0 397
rect -88 285 0 351
rect -88 239 -75 285
rect -29 239 0 285
rect -88 172 0 239
rect -88 126 -75 172
rect -29 126 0 172
rect -88 59 0 126
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 509 224 522
rect 120 463 149 509
rect 195 463 224 509
rect 120 397 224 463
rect 120 351 149 397
rect 195 351 224 397
rect 120 285 224 351
rect 120 239 149 285
rect 195 239 224 285
rect 120 172 224 239
rect 120 126 149 172
rect 195 126 224 172
rect 120 59 224 126
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 509 432 522
rect 344 463 373 509
rect 419 463 432 509
rect 344 397 432 463
rect 344 351 373 397
rect 419 351 432 397
rect 344 285 432 351
rect 344 239 373 285
rect 419 239 432 285
rect 344 172 432 239
rect 344 126 373 172
rect 419 126 432 172
rect 344 59 432 126
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvndiffc >>
rect -75 463 -29 509
rect -75 351 -29 397
rect -75 239 -29 285
rect -75 126 -29 172
rect -75 13 -29 59
rect 149 463 195 509
rect 149 351 195 397
rect 149 239 195 285
rect 149 126 195 172
rect 149 13 195 59
rect 373 463 419 509
rect 373 351 419 397
rect 373 239 419 285
rect 373 126 419 172
rect 373 13 419 59
<< polysilicon >>
rect 0 522 120 566
rect 224 522 344 566
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 509 -29 522
rect -75 397 -29 463
rect -75 285 -29 351
rect -75 172 -29 239
rect -75 59 -29 126
rect -75 0 -29 13
rect 149 509 195 522
rect 149 397 195 463
rect 149 285 195 351
rect 149 172 195 239
rect 149 59 195 126
rect 149 0 195 13
rect 373 509 419 522
rect 373 397 419 463
rect 373 285 419 351
rect 373 172 419 239
rect 373 59 419 126
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 261 -52 261 0 FreeSans 200 0 0 0 S
flabel metal1 s 396 261 396 261 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 261 172 261 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 147904
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 145666
<< end >>
