magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 364
rect 224 0 344 364
<< mvndiff >>
rect -88 351 0 364
rect -88 305 -75 351
rect -29 305 0 351
rect -88 205 0 305
rect -88 159 -75 205
rect -29 159 0 205
rect -88 59 0 159
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 351 224 364
rect 120 305 149 351
rect 195 305 224 351
rect 120 205 224 305
rect 120 159 149 205
rect 195 159 224 205
rect 120 59 224 159
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 351 432 364
rect 344 305 373 351
rect 419 305 432 351
rect 344 205 432 305
rect 344 159 373 205
rect 419 159 432 205
rect 344 59 432 159
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvndiffc >>
rect -75 305 -29 351
rect -75 159 -29 205
rect -75 13 -29 59
rect 149 305 195 351
rect 149 159 195 205
rect 149 13 195 59
rect 373 305 419 351
rect 373 159 419 205
rect 373 13 419 59
<< polysilicon >>
rect 0 364 120 408
rect 224 364 344 408
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 351 -29 364
rect -75 205 -29 305
rect -75 59 -29 159
rect -75 0 -29 13
rect 149 351 195 364
rect 149 205 195 305
rect 149 59 195 159
rect 149 0 195 13
rect 373 351 419 364
rect 373 205 419 305
rect 373 59 419 159
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 182 -52 182 0 FreeSans 200 0 0 0 S
flabel metal1 s 396 182 396 182 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 182 172 182 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 2006
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 152
<< end >>
