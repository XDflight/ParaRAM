magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 454 88 527
rect 193 454 312 527
rect -31 -73 88 -1
rect 193 -73 312 -1
use nmos_5p04310590878139_256x8m81  nmos_5p04310590878139_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 432 498
<< properties >>
string GDS_END 1094960
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1094582
<< end >>
