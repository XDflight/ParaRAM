magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -546 -142 344 3179
<< polysilicon >>
rect -31 3039 88 3111
rect -31 -74 88 -1
use pmos_5p04310590548771_128x8m81  pmos_5p04310590548771_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 3160
<< properties >>
string GDS_END 214332
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 213954
<< end >>
