magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 1028
<< mvpmos >>
rect 0 0 120 908
rect 224 0 344 908
<< mvpdiff >>
rect -88 895 0 908
rect -88 849 -75 895
rect -29 849 0 895
rect -88 791 0 849
rect -88 745 -75 791
rect -29 745 0 791
rect -88 687 0 745
rect -88 641 -75 687
rect -29 641 0 687
rect -88 583 0 641
rect -88 537 -75 583
rect -29 537 0 583
rect -88 479 0 537
rect -88 433 -75 479
rect -29 433 0 479
rect -88 374 0 433
rect -88 328 -75 374
rect -29 328 0 374
rect -88 269 0 328
rect -88 223 -75 269
rect -29 223 0 269
rect -88 164 0 223
rect -88 118 -75 164
rect -29 118 0 164
rect -88 59 0 118
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 895 224 908
rect 120 849 149 895
rect 195 849 224 895
rect 120 791 224 849
rect 120 745 149 791
rect 195 745 224 791
rect 120 687 224 745
rect 120 641 149 687
rect 195 641 224 687
rect 120 583 224 641
rect 120 537 149 583
rect 195 537 224 583
rect 120 479 224 537
rect 120 433 149 479
rect 195 433 224 479
rect 120 374 224 433
rect 120 328 149 374
rect 195 328 224 374
rect 120 269 224 328
rect 120 223 149 269
rect 195 223 224 269
rect 120 164 224 223
rect 120 118 149 164
rect 195 118 224 164
rect 120 59 224 118
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 895 432 908
rect 344 849 373 895
rect 419 849 432 895
rect 344 791 432 849
rect 344 745 373 791
rect 419 745 432 791
rect 344 687 432 745
rect 344 641 373 687
rect 419 641 432 687
rect 344 583 432 641
rect 344 537 373 583
rect 419 537 432 583
rect 344 479 432 537
rect 344 433 373 479
rect 419 433 432 479
rect 344 374 432 433
rect 344 328 373 374
rect 419 328 432 374
rect 344 269 432 328
rect 344 223 373 269
rect 419 223 432 269
rect 344 164 432 223
rect 344 118 373 164
rect 419 118 432 164
rect 344 59 432 118
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 849 -29 895
rect -75 745 -29 791
rect -75 641 -29 687
rect -75 537 -29 583
rect -75 433 -29 479
rect -75 328 -29 374
rect -75 223 -29 269
rect -75 118 -29 164
rect -75 13 -29 59
rect 149 849 195 895
rect 149 745 195 791
rect 149 641 195 687
rect 149 537 195 583
rect 149 433 195 479
rect 149 328 195 374
rect 149 223 195 269
rect 149 118 195 164
rect 149 13 195 59
rect 373 849 419 895
rect 373 745 419 791
rect 373 641 419 687
rect 373 537 419 583
rect 373 433 419 479
rect 373 328 419 374
rect 373 223 419 269
rect 373 118 419 164
rect 373 13 419 59
<< polysilicon >>
rect 0 908 120 952
rect 224 908 344 952
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 895 -29 908
rect -75 791 -29 849
rect -75 687 -29 745
rect -75 583 -29 641
rect -75 479 -29 537
rect -75 374 -29 433
rect -75 269 -29 328
rect -75 164 -29 223
rect -75 59 -29 118
rect -75 0 -29 13
rect 149 895 195 908
rect 149 791 195 849
rect 149 687 195 745
rect 149 583 195 641
rect 149 479 195 537
rect 149 374 195 433
rect 149 269 195 328
rect 149 164 195 223
rect 149 59 195 118
rect 149 0 195 13
rect 373 895 419 908
rect 373 791 419 849
rect 373 687 419 745
rect 373 583 419 641
rect 373 479 419 537
rect 373 374 419 433
rect 373 269 419 328
rect 373 164 419 223
rect 373 59 419 118
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 454 -52 454 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 454 396 454 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 454 172 454 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 12630
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 9560
<< end >>
