magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -1029 23 1029 42
rect -1029 -23 -1010 23
rect 1010 -23 1029 23
rect -1029 -42 1029 -23
<< polycontact >>
rect -1010 -23 1010 23
<< metal1 >>
rect -1021 23 1021 34
rect -1021 -23 -1010 23
rect 1010 -23 1021 23
rect -1021 -34 1021 -23
<< properties >>
string GDS_END 1037810
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1036270
<< end >>
