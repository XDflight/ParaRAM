magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -1975 39 1975 58
rect -1975 -7 -1762 39
rect -1716 -7 -1604 39
rect -1558 -7 -1446 39
rect -1400 -7 -1288 39
rect -1242 -7 -1130 39
rect -1084 -7 -972 39
rect -926 -7 -814 39
rect -768 -7 -656 39
rect -610 -7 -497 39
rect -451 -7 -339 39
rect -293 -7 -181 39
rect -135 -7 -23 39
rect 23 -7 135 39
rect 181 -7 293 39
rect 339 -7 451 39
rect 497 -7 610 39
rect 656 -7 768 39
rect 814 -7 926 39
rect 972 -7 1084 39
rect 1130 -7 1242 39
rect 1288 -7 1400 39
rect 1446 -7 1558 39
rect 1604 -7 1716 39
rect 1762 -7 1874 39
rect 1920 -7 1975 39
rect -1975 -26 1975 -7
<< psubdiffcont >>
rect -1762 -7 -1716 39
rect -1604 -7 -1558 39
rect -1446 -7 -1400 39
rect -1288 -7 -1242 39
rect -1130 -7 -1084 39
rect -972 -7 -926 39
rect -814 -7 -768 39
rect -656 -7 -610 39
rect -497 -7 -451 39
rect -339 -7 -293 39
rect -181 -7 -135 39
rect -23 -7 23 39
rect 135 -7 181 39
rect 293 -7 339 39
rect 451 -7 497 39
rect 610 -7 656 39
rect 768 -7 814 39
rect 926 -7 972 39
rect 1084 -7 1130 39
rect 1242 -7 1288 39
rect 1400 -7 1446 39
rect 1558 -7 1604 39
rect 1716 -7 1762 39
rect 1874 -7 1920 39
<< metal1 >>
rect -1955 39 1955 50
rect -1955 -7 -1762 39
rect -1716 -7 -1604 39
rect -1558 -7 -1446 39
rect -1400 -7 -1288 39
rect -1242 -7 -1130 39
rect -1084 -7 -972 39
rect -926 -7 -814 39
rect -768 -7 -656 39
rect -610 -7 -497 39
rect -451 -7 -339 39
rect -293 -7 -181 39
rect -135 -7 -23 39
rect 23 -7 135 39
rect 181 -7 293 39
rect 339 -7 451 39
rect 497 -7 610 39
rect 656 -7 768 39
rect 814 -7 926 39
rect 972 -7 1084 39
rect 1130 -7 1242 39
rect 1288 -7 1400 39
rect 1446 -7 1558 39
rect 1604 -7 1716 39
rect 1762 -7 1874 39
rect 1920 -7 1955 39
rect -1955 -18 1955 -7
<< properties >>
string GDS_END 380460
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 378728
<< end >>
