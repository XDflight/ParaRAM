magic
tech gf180mcuC
magscale 1 5
timestamp 1667831717
<< obsm1 >>
rect 672 1538 299320 299809
<< metal2 >>
rect 4900 299760 5012 300480
rect 13188 299760 13300 300480
rect 21476 299760 21588 300480
rect 29764 299760 29876 300480
rect 38052 299760 38164 300480
rect 46340 299760 46452 300480
rect 54628 299760 54740 300480
rect 62916 299760 63028 300480
rect 71204 299760 71316 300480
rect 79492 299760 79604 300480
rect 87780 299760 87892 300480
rect 96068 299760 96180 300480
rect 104356 299760 104468 300480
rect 112644 299760 112756 300480
rect 120932 299760 121044 300480
rect 129220 299760 129332 300480
rect 137508 299760 137620 300480
rect 145796 299760 145908 300480
rect 154084 299760 154196 300480
rect 162372 299760 162484 300480
rect 170660 299760 170772 300480
rect 178948 299760 179060 300480
rect 187236 299760 187348 300480
rect 195524 299760 195636 300480
rect 203812 299760 203924 300480
rect 212100 299760 212212 300480
rect 220388 299760 220500 300480
rect 228676 299760 228788 300480
rect 236964 299760 237076 300480
rect 245252 299760 245364 300480
rect 253540 299760 253652 300480
rect 261828 299760 261940 300480
rect 270116 299760 270228 300480
rect 278404 299760 278516 300480
rect 286692 299760 286804 300480
rect 294980 299760 295092 300480
rect 11900 -480 12012 240
rect 12460 -480 12572 240
rect 13020 -480 13132 240
rect 13580 -480 13692 240
rect 14140 -480 14252 240
rect 14700 -480 14812 240
rect 15260 -480 15372 240
rect 15820 -480 15932 240
rect 16380 -480 16492 240
rect 16940 -480 17052 240
rect 17500 -480 17612 240
rect 18060 -480 18172 240
rect 18620 -480 18732 240
rect 19180 -480 19292 240
rect 19740 -480 19852 240
rect 20300 -480 20412 240
rect 20860 -480 20972 240
rect 21420 -480 21532 240
rect 21980 -480 22092 240
rect 22540 -480 22652 240
rect 23100 -480 23212 240
rect 23660 -480 23772 240
rect 24220 -480 24332 240
rect 24780 -480 24892 240
rect 25340 -480 25452 240
rect 25900 -480 26012 240
rect 26460 -480 26572 240
rect 27020 -480 27132 240
rect 27580 -480 27692 240
rect 28140 -480 28252 240
rect 28700 -480 28812 240
rect 29260 -480 29372 240
rect 29820 -480 29932 240
rect 30380 -480 30492 240
rect 30940 -480 31052 240
rect 31500 -480 31612 240
rect 32060 -480 32172 240
rect 32620 -480 32732 240
rect 33180 -480 33292 240
rect 33740 -480 33852 240
rect 34300 -480 34412 240
rect 34860 -480 34972 240
rect 35420 -480 35532 240
rect 35980 -480 36092 240
rect 36540 -480 36652 240
rect 37100 -480 37212 240
rect 37660 -480 37772 240
rect 38220 -480 38332 240
rect 38780 -480 38892 240
rect 39340 -480 39452 240
rect 39900 -480 40012 240
rect 40460 -480 40572 240
rect 41020 -480 41132 240
rect 41580 -480 41692 240
rect 42140 -480 42252 240
rect 42700 -480 42812 240
rect 43260 -480 43372 240
rect 43820 -480 43932 240
rect 44380 -480 44492 240
rect 44940 -480 45052 240
rect 45500 -480 45612 240
rect 46060 -480 46172 240
rect 46620 -480 46732 240
rect 47180 -480 47292 240
rect 47740 -480 47852 240
rect 48300 -480 48412 240
rect 48860 -480 48972 240
rect 49420 -480 49532 240
rect 49980 -480 50092 240
rect 50540 -480 50652 240
rect 51100 -480 51212 240
rect 51660 -480 51772 240
rect 52220 -480 52332 240
rect 52780 -480 52892 240
rect 53340 -480 53452 240
rect 53900 -480 54012 240
rect 54460 -480 54572 240
rect 55020 -480 55132 240
rect 55580 -480 55692 240
rect 56140 -480 56252 240
rect 56700 -480 56812 240
rect 57260 -480 57372 240
rect 57820 -480 57932 240
rect 58380 -480 58492 240
rect 58940 -480 59052 240
rect 59500 -480 59612 240
rect 60060 -480 60172 240
rect 60620 -480 60732 240
rect 61180 -480 61292 240
rect 61740 -480 61852 240
rect 62300 -480 62412 240
rect 62860 -480 62972 240
rect 63420 -480 63532 240
rect 63980 -480 64092 240
rect 64540 -480 64652 240
rect 65100 -480 65212 240
rect 65660 -480 65772 240
rect 66220 -480 66332 240
rect 66780 -480 66892 240
rect 67340 -480 67452 240
rect 67900 -480 68012 240
rect 68460 -480 68572 240
rect 69020 -480 69132 240
rect 69580 -480 69692 240
rect 70140 -480 70252 240
rect 70700 -480 70812 240
rect 71260 -480 71372 240
rect 71820 -480 71932 240
rect 72380 -480 72492 240
rect 72940 -480 73052 240
rect 73500 -480 73612 240
rect 74060 -480 74172 240
rect 74620 -480 74732 240
rect 75180 -480 75292 240
rect 75740 -480 75852 240
rect 76300 -480 76412 240
rect 76860 -480 76972 240
rect 77420 -480 77532 240
rect 77980 -480 78092 240
rect 78540 -480 78652 240
rect 79100 -480 79212 240
rect 79660 -480 79772 240
rect 80220 -480 80332 240
rect 80780 -480 80892 240
rect 81340 -480 81452 240
rect 81900 -480 82012 240
rect 82460 -480 82572 240
rect 83020 -480 83132 240
rect 83580 -480 83692 240
rect 84140 -480 84252 240
rect 84700 -480 84812 240
rect 85260 -480 85372 240
rect 85820 -480 85932 240
rect 86380 -480 86492 240
rect 86940 -480 87052 240
rect 87500 -480 87612 240
rect 88060 -480 88172 240
rect 88620 -480 88732 240
rect 89180 -480 89292 240
rect 89740 -480 89852 240
rect 90300 -480 90412 240
rect 90860 -480 90972 240
rect 91420 -480 91532 240
rect 91980 -480 92092 240
rect 92540 -480 92652 240
rect 93100 -480 93212 240
rect 93660 -480 93772 240
rect 94220 -480 94332 240
rect 94780 -480 94892 240
rect 95340 -480 95452 240
rect 95900 -480 96012 240
rect 96460 -480 96572 240
rect 97020 -480 97132 240
rect 97580 -480 97692 240
rect 98140 -480 98252 240
rect 98700 -480 98812 240
rect 99260 -480 99372 240
rect 99820 -480 99932 240
rect 100380 -480 100492 240
rect 100940 -480 101052 240
rect 101500 -480 101612 240
rect 102060 -480 102172 240
rect 102620 -480 102732 240
rect 103180 -480 103292 240
rect 103740 -480 103852 240
rect 104300 -480 104412 240
rect 104860 -480 104972 240
rect 105420 -480 105532 240
rect 105980 -480 106092 240
rect 106540 -480 106652 240
rect 107100 -480 107212 240
rect 107660 -480 107772 240
rect 108220 -480 108332 240
rect 108780 -480 108892 240
rect 109340 -480 109452 240
rect 109900 -480 110012 240
rect 110460 -480 110572 240
rect 111020 -480 111132 240
rect 111580 -480 111692 240
rect 112140 -480 112252 240
rect 112700 -480 112812 240
rect 113260 -480 113372 240
rect 113820 -480 113932 240
rect 114380 -480 114492 240
rect 114940 -480 115052 240
rect 115500 -480 115612 240
rect 116060 -480 116172 240
rect 116620 -480 116732 240
rect 117180 -480 117292 240
rect 117740 -480 117852 240
rect 118300 -480 118412 240
rect 118860 -480 118972 240
rect 119420 -480 119532 240
rect 119980 -480 120092 240
rect 120540 -480 120652 240
rect 121100 -480 121212 240
rect 121660 -480 121772 240
rect 122220 -480 122332 240
rect 122780 -480 122892 240
rect 123340 -480 123452 240
rect 123900 -480 124012 240
rect 124460 -480 124572 240
rect 125020 -480 125132 240
rect 125580 -480 125692 240
rect 126140 -480 126252 240
rect 126700 -480 126812 240
rect 127260 -480 127372 240
rect 127820 -480 127932 240
rect 128380 -480 128492 240
rect 128940 -480 129052 240
rect 129500 -480 129612 240
rect 130060 -480 130172 240
rect 130620 -480 130732 240
rect 131180 -480 131292 240
rect 131740 -480 131852 240
rect 132300 -480 132412 240
rect 132860 -480 132972 240
rect 133420 -480 133532 240
rect 133980 -480 134092 240
rect 134540 -480 134652 240
rect 135100 -480 135212 240
rect 135660 -480 135772 240
rect 136220 -480 136332 240
rect 136780 -480 136892 240
rect 137340 -480 137452 240
rect 137900 -480 138012 240
rect 138460 -480 138572 240
rect 139020 -480 139132 240
rect 139580 -480 139692 240
rect 140140 -480 140252 240
rect 140700 -480 140812 240
rect 141260 -480 141372 240
rect 141820 -480 141932 240
rect 142380 -480 142492 240
rect 142940 -480 143052 240
rect 143500 -480 143612 240
rect 144060 -480 144172 240
rect 144620 -480 144732 240
rect 145180 -480 145292 240
rect 145740 -480 145852 240
rect 146300 -480 146412 240
rect 146860 -480 146972 240
rect 147420 -480 147532 240
rect 147980 -480 148092 240
rect 148540 -480 148652 240
rect 149100 -480 149212 240
rect 149660 -480 149772 240
rect 150220 -480 150332 240
rect 150780 -480 150892 240
rect 151340 -480 151452 240
rect 151900 -480 152012 240
rect 152460 -480 152572 240
rect 153020 -480 153132 240
rect 153580 -480 153692 240
rect 154140 -480 154252 240
rect 154700 -480 154812 240
rect 155260 -480 155372 240
rect 155820 -480 155932 240
rect 156380 -480 156492 240
rect 156940 -480 157052 240
rect 157500 -480 157612 240
rect 158060 -480 158172 240
rect 158620 -480 158732 240
rect 159180 -480 159292 240
rect 159740 -480 159852 240
rect 160300 -480 160412 240
rect 160860 -480 160972 240
rect 161420 -480 161532 240
rect 161980 -480 162092 240
rect 162540 -480 162652 240
rect 163100 -480 163212 240
rect 163660 -480 163772 240
rect 164220 -480 164332 240
rect 164780 -480 164892 240
rect 165340 -480 165452 240
rect 165900 -480 166012 240
rect 166460 -480 166572 240
rect 167020 -480 167132 240
rect 167580 -480 167692 240
rect 168140 -480 168252 240
rect 168700 -480 168812 240
rect 169260 -480 169372 240
rect 169820 -480 169932 240
rect 170380 -480 170492 240
rect 170940 -480 171052 240
rect 171500 -480 171612 240
rect 172060 -480 172172 240
rect 172620 -480 172732 240
rect 173180 -480 173292 240
rect 173740 -480 173852 240
rect 174300 -480 174412 240
rect 174860 -480 174972 240
rect 175420 -480 175532 240
rect 175980 -480 176092 240
rect 176540 -480 176652 240
rect 177100 -480 177212 240
rect 177660 -480 177772 240
rect 178220 -480 178332 240
rect 178780 -480 178892 240
rect 179340 -480 179452 240
rect 179900 -480 180012 240
rect 180460 -480 180572 240
rect 181020 -480 181132 240
rect 181580 -480 181692 240
rect 182140 -480 182252 240
rect 182700 -480 182812 240
rect 183260 -480 183372 240
rect 183820 -480 183932 240
rect 184380 -480 184492 240
rect 184940 -480 185052 240
rect 185500 -480 185612 240
rect 186060 -480 186172 240
rect 186620 -480 186732 240
rect 187180 -480 187292 240
rect 187740 -480 187852 240
rect 188300 -480 188412 240
rect 188860 -480 188972 240
rect 189420 -480 189532 240
rect 189980 -480 190092 240
rect 190540 -480 190652 240
rect 191100 -480 191212 240
rect 191660 -480 191772 240
rect 192220 -480 192332 240
rect 192780 -480 192892 240
rect 193340 -480 193452 240
rect 193900 -480 194012 240
rect 194460 -480 194572 240
rect 195020 -480 195132 240
rect 195580 -480 195692 240
rect 196140 -480 196252 240
rect 196700 -480 196812 240
rect 197260 -480 197372 240
rect 197820 -480 197932 240
rect 198380 -480 198492 240
rect 198940 -480 199052 240
rect 199500 -480 199612 240
rect 200060 -480 200172 240
rect 200620 -480 200732 240
rect 201180 -480 201292 240
rect 201740 -480 201852 240
rect 202300 -480 202412 240
rect 202860 -480 202972 240
rect 203420 -480 203532 240
rect 203980 -480 204092 240
rect 204540 -480 204652 240
rect 205100 -480 205212 240
rect 205660 -480 205772 240
rect 206220 -480 206332 240
rect 206780 -480 206892 240
rect 207340 -480 207452 240
rect 207900 -480 208012 240
rect 208460 -480 208572 240
rect 209020 -480 209132 240
rect 209580 -480 209692 240
rect 210140 -480 210252 240
rect 210700 -480 210812 240
rect 211260 -480 211372 240
rect 211820 -480 211932 240
rect 212380 -480 212492 240
rect 212940 -480 213052 240
rect 213500 -480 213612 240
rect 214060 -480 214172 240
rect 214620 -480 214732 240
rect 215180 -480 215292 240
rect 215740 -480 215852 240
rect 216300 -480 216412 240
rect 216860 -480 216972 240
rect 217420 -480 217532 240
rect 217980 -480 218092 240
rect 218540 -480 218652 240
rect 219100 -480 219212 240
rect 219660 -480 219772 240
rect 220220 -480 220332 240
rect 220780 -480 220892 240
rect 221340 -480 221452 240
rect 221900 -480 222012 240
rect 222460 -480 222572 240
rect 223020 -480 223132 240
rect 223580 -480 223692 240
rect 224140 -480 224252 240
rect 224700 -480 224812 240
rect 225260 -480 225372 240
rect 225820 -480 225932 240
rect 226380 -480 226492 240
rect 226940 -480 227052 240
rect 227500 -480 227612 240
rect 228060 -480 228172 240
rect 228620 -480 228732 240
rect 229180 -480 229292 240
rect 229740 -480 229852 240
rect 230300 -480 230412 240
rect 230860 -480 230972 240
rect 231420 -480 231532 240
rect 231980 -480 232092 240
rect 232540 -480 232652 240
rect 233100 -480 233212 240
rect 233660 -480 233772 240
rect 234220 -480 234332 240
rect 234780 -480 234892 240
rect 235340 -480 235452 240
rect 235900 -480 236012 240
rect 236460 -480 236572 240
rect 237020 -480 237132 240
rect 237580 -480 237692 240
rect 238140 -480 238252 240
rect 238700 -480 238812 240
rect 239260 -480 239372 240
rect 239820 -480 239932 240
rect 240380 -480 240492 240
rect 240940 -480 241052 240
rect 241500 -480 241612 240
rect 242060 -480 242172 240
rect 242620 -480 242732 240
rect 243180 -480 243292 240
rect 243740 -480 243852 240
rect 244300 -480 244412 240
rect 244860 -480 244972 240
rect 245420 -480 245532 240
rect 245980 -480 246092 240
rect 246540 -480 246652 240
rect 247100 -480 247212 240
rect 247660 -480 247772 240
rect 248220 -480 248332 240
rect 248780 -480 248892 240
rect 249340 -480 249452 240
rect 249900 -480 250012 240
rect 250460 -480 250572 240
rect 251020 -480 251132 240
rect 251580 -480 251692 240
rect 252140 -480 252252 240
rect 252700 -480 252812 240
rect 253260 -480 253372 240
rect 253820 -480 253932 240
rect 254380 -480 254492 240
rect 254940 -480 255052 240
rect 255500 -480 255612 240
rect 256060 -480 256172 240
rect 256620 -480 256732 240
rect 257180 -480 257292 240
rect 257740 -480 257852 240
rect 258300 -480 258412 240
rect 258860 -480 258972 240
rect 259420 -480 259532 240
rect 259980 -480 260092 240
rect 260540 -480 260652 240
rect 261100 -480 261212 240
rect 261660 -480 261772 240
rect 262220 -480 262332 240
rect 262780 -480 262892 240
rect 263340 -480 263452 240
rect 263900 -480 264012 240
rect 264460 -480 264572 240
rect 265020 -480 265132 240
rect 265580 -480 265692 240
rect 266140 -480 266252 240
rect 266700 -480 266812 240
rect 267260 -480 267372 240
rect 267820 -480 267932 240
rect 268380 -480 268492 240
rect 268940 -480 269052 240
rect 269500 -480 269612 240
rect 270060 -480 270172 240
rect 270620 -480 270732 240
rect 271180 -480 271292 240
rect 271740 -480 271852 240
rect 272300 -480 272412 240
rect 272860 -480 272972 240
rect 273420 -480 273532 240
rect 273980 -480 274092 240
rect 274540 -480 274652 240
rect 275100 -480 275212 240
rect 275660 -480 275772 240
rect 276220 -480 276332 240
rect 276780 -480 276892 240
rect 277340 -480 277452 240
rect 277900 -480 278012 240
rect 278460 -480 278572 240
rect 279020 -480 279132 240
rect 279580 -480 279692 240
rect 280140 -480 280252 240
rect 280700 -480 280812 240
rect 281260 -480 281372 240
rect 281820 -480 281932 240
rect 282380 -480 282492 240
rect 282940 -480 283052 240
rect 283500 -480 283612 240
rect 284060 -480 284172 240
rect 284620 -480 284732 240
rect 285180 -480 285292 240
rect 285740 -480 285852 240
rect 286300 -480 286412 240
rect 286860 -480 286972 240
rect 287420 -480 287532 240
rect 287980 -480 288092 240
<< obsm2 >>
rect 910 299730 4870 299983
rect 5042 299730 13158 299983
rect 13330 299730 21446 299983
rect 21618 299730 29734 299983
rect 29906 299730 38022 299983
rect 38194 299730 46310 299983
rect 46482 299730 54598 299983
rect 54770 299730 62886 299983
rect 63058 299730 71174 299983
rect 71346 299730 79462 299983
rect 79634 299730 87750 299983
rect 87922 299730 96038 299983
rect 96210 299730 104326 299983
rect 104498 299730 112614 299983
rect 112786 299730 120902 299983
rect 121074 299730 129190 299983
rect 129362 299730 137478 299983
rect 137650 299730 145766 299983
rect 145938 299730 154054 299983
rect 154226 299730 162342 299983
rect 162514 299730 170630 299983
rect 170802 299730 178918 299983
rect 179090 299730 187206 299983
rect 187378 299730 195494 299983
rect 195666 299730 203782 299983
rect 203954 299730 212070 299983
rect 212242 299730 220358 299983
rect 220530 299730 228646 299983
rect 228818 299730 236934 299983
rect 237106 299730 245222 299983
rect 245394 299730 253510 299983
rect 253682 299730 261798 299983
rect 261970 299730 270086 299983
rect 270258 299730 278374 299983
rect 278546 299730 286662 299983
rect 286834 299730 294950 299983
rect 295122 299730 299082 299983
rect 910 270 299082 299730
rect 910 182 11870 270
rect 12042 182 12430 270
rect 12602 182 12990 270
rect 13162 182 13550 270
rect 13722 182 14110 270
rect 14282 182 14670 270
rect 14842 182 15230 270
rect 15402 182 15790 270
rect 15962 182 16350 270
rect 16522 182 16910 270
rect 17082 182 17470 270
rect 17642 182 18030 270
rect 18202 182 18590 270
rect 18762 182 19150 270
rect 19322 182 19710 270
rect 19882 182 20270 270
rect 20442 182 20830 270
rect 21002 182 21390 270
rect 21562 182 21950 270
rect 22122 182 22510 270
rect 22682 182 23070 270
rect 23242 182 23630 270
rect 23802 182 24190 270
rect 24362 182 24750 270
rect 24922 182 25310 270
rect 25482 182 25870 270
rect 26042 182 26430 270
rect 26602 182 26990 270
rect 27162 182 27550 270
rect 27722 182 28110 270
rect 28282 182 28670 270
rect 28842 182 29230 270
rect 29402 182 29790 270
rect 29962 182 30350 270
rect 30522 182 30910 270
rect 31082 182 31470 270
rect 31642 182 32030 270
rect 32202 182 32590 270
rect 32762 182 33150 270
rect 33322 182 33710 270
rect 33882 182 34270 270
rect 34442 182 34830 270
rect 35002 182 35390 270
rect 35562 182 35950 270
rect 36122 182 36510 270
rect 36682 182 37070 270
rect 37242 182 37630 270
rect 37802 182 38190 270
rect 38362 182 38750 270
rect 38922 182 39310 270
rect 39482 182 39870 270
rect 40042 182 40430 270
rect 40602 182 40990 270
rect 41162 182 41550 270
rect 41722 182 42110 270
rect 42282 182 42670 270
rect 42842 182 43230 270
rect 43402 182 43790 270
rect 43962 182 44350 270
rect 44522 182 44910 270
rect 45082 182 45470 270
rect 45642 182 46030 270
rect 46202 182 46590 270
rect 46762 182 47150 270
rect 47322 182 47710 270
rect 47882 182 48270 270
rect 48442 182 48830 270
rect 49002 182 49390 270
rect 49562 182 49950 270
rect 50122 182 50510 270
rect 50682 182 51070 270
rect 51242 182 51630 270
rect 51802 182 52190 270
rect 52362 182 52750 270
rect 52922 182 53310 270
rect 53482 182 53870 270
rect 54042 182 54430 270
rect 54602 182 54990 270
rect 55162 182 55550 270
rect 55722 182 56110 270
rect 56282 182 56670 270
rect 56842 182 57230 270
rect 57402 182 57790 270
rect 57962 182 58350 270
rect 58522 182 58910 270
rect 59082 182 59470 270
rect 59642 182 60030 270
rect 60202 182 60590 270
rect 60762 182 61150 270
rect 61322 182 61710 270
rect 61882 182 62270 270
rect 62442 182 62830 270
rect 63002 182 63390 270
rect 63562 182 63950 270
rect 64122 182 64510 270
rect 64682 182 65070 270
rect 65242 182 65630 270
rect 65802 182 66190 270
rect 66362 182 66750 270
rect 66922 182 67310 270
rect 67482 182 67870 270
rect 68042 182 68430 270
rect 68602 182 68990 270
rect 69162 182 69550 270
rect 69722 182 70110 270
rect 70282 182 70670 270
rect 70842 182 71230 270
rect 71402 182 71790 270
rect 71962 182 72350 270
rect 72522 182 72910 270
rect 73082 182 73470 270
rect 73642 182 74030 270
rect 74202 182 74590 270
rect 74762 182 75150 270
rect 75322 182 75710 270
rect 75882 182 76270 270
rect 76442 182 76830 270
rect 77002 182 77390 270
rect 77562 182 77950 270
rect 78122 182 78510 270
rect 78682 182 79070 270
rect 79242 182 79630 270
rect 79802 182 80190 270
rect 80362 182 80750 270
rect 80922 182 81310 270
rect 81482 182 81870 270
rect 82042 182 82430 270
rect 82602 182 82990 270
rect 83162 182 83550 270
rect 83722 182 84110 270
rect 84282 182 84670 270
rect 84842 182 85230 270
rect 85402 182 85790 270
rect 85962 182 86350 270
rect 86522 182 86910 270
rect 87082 182 87470 270
rect 87642 182 88030 270
rect 88202 182 88590 270
rect 88762 182 89150 270
rect 89322 182 89710 270
rect 89882 182 90270 270
rect 90442 182 90830 270
rect 91002 182 91390 270
rect 91562 182 91950 270
rect 92122 182 92510 270
rect 92682 182 93070 270
rect 93242 182 93630 270
rect 93802 182 94190 270
rect 94362 182 94750 270
rect 94922 182 95310 270
rect 95482 182 95870 270
rect 96042 182 96430 270
rect 96602 182 96990 270
rect 97162 182 97550 270
rect 97722 182 98110 270
rect 98282 182 98670 270
rect 98842 182 99230 270
rect 99402 182 99790 270
rect 99962 182 100350 270
rect 100522 182 100910 270
rect 101082 182 101470 270
rect 101642 182 102030 270
rect 102202 182 102590 270
rect 102762 182 103150 270
rect 103322 182 103710 270
rect 103882 182 104270 270
rect 104442 182 104830 270
rect 105002 182 105390 270
rect 105562 182 105950 270
rect 106122 182 106510 270
rect 106682 182 107070 270
rect 107242 182 107630 270
rect 107802 182 108190 270
rect 108362 182 108750 270
rect 108922 182 109310 270
rect 109482 182 109870 270
rect 110042 182 110430 270
rect 110602 182 110990 270
rect 111162 182 111550 270
rect 111722 182 112110 270
rect 112282 182 112670 270
rect 112842 182 113230 270
rect 113402 182 113790 270
rect 113962 182 114350 270
rect 114522 182 114910 270
rect 115082 182 115470 270
rect 115642 182 116030 270
rect 116202 182 116590 270
rect 116762 182 117150 270
rect 117322 182 117710 270
rect 117882 182 118270 270
rect 118442 182 118830 270
rect 119002 182 119390 270
rect 119562 182 119950 270
rect 120122 182 120510 270
rect 120682 182 121070 270
rect 121242 182 121630 270
rect 121802 182 122190 270
rect 122362 182 122750 270
rect 122922 182 123310 270
rect 123482 182 123870 270
rect 124042 182 124430 270
rect 124602 182 124990 270
rect 125162 182 125550 270
rect 125722 182 126110 270
rect 126282 182 126670 270
rect 126842 182 127230 270
rect 127402 182 127790 270
rect 127962 182 128350 270
rect 128522 182 128910 270
rect 129082 182 129470 270
rect 129642 182 130030 270
rect 130202 182 130590 270
rect 130762 182 131150 270
rect 131322 182 131710 270
rect 131882 182 132270 270
rect 132442 182 132830 270
rect 133002 182 133390 270
rect 133562 182 133950 270
rect 134122 182 134510 270
rect 134682 182 135070 270
rect 135242 182 135630 270
rect 135802 182 136190 270
rect 136362 182 136750 270
rect 136922 182 137310 270
rect 137482 182 137870 270
rect 138042 182 138430 270
rect 138602 182 138990 270
rect 139162 182 139550 270
rect 139722 182 140110 270
rect 140282 182 140670 270
rect 140842 182 141230 270
rect 141402 182 141790 270
rect 141962 182 142350 270
rect 142522 182 142910 270
rect 143082 182 143470 270
rect 143642 182 144030 270
rect 144202 182 144590 270
rect 144762 182 145150 270
rect 145322 182 145710 270
rect 145882 182 146270 270
rect 146442 182 146830 270
rect 147002 182 147390 270
rect 147562 182 147950 270
rect 148122 182 148510 270
rect 148682 182 149070 270
rect 149242 182 149630 270
rect 149802 182 150190 270
rect 150362 182 150750 270
rect 150922 182 151310 270
rect 151482 182 151870 270
rect 152042 182 152430 270
rect 152602 182 152990 270
rect 153162 182 153550 270
rect 153722 182 154110 270
rect 154282 182 154670 270
rect 154842 182 155230 270
rect 155402 182 155790 270
rect 155962 182 156350 270
rect 156522 182 156910 270
rect 157082 182 157470 270
rect 157642 182 158030 270
rect 158202 182 158590 270
rect 158762 182 159150 270
rect 159322 182 159710 270
rect 159882 182 160270 270
rect 160442 182 160830 270
rect 161002 182 161390 270
rect 161562 182 161950 270
rect 162122 182 162510 270
rect 162682 182 163070 270
rect 163242 182 163630 270
rect 163802 182 164190 270
rect 164362 182 164750 270
rect 164922 182 165310 270
rect 165482 182 165870 270
rect 166042 182 166430 270
rect 166602 182 166990 270
rect 167162 182 167550 270
rect 167722 182 168110 270
rect 168282 182 168670 270
rect 168842 182 169230 270
rect 169402 182 169790 270
rect 169962 182 170350 270
rect 170522 182 170910 270
rect 171082 182 171470 270
rect 171642 182 172030 270
rect 172202 182 172590 270
rect 172762 182 173150 270
rect 173322 182 173710 270
rect 173882 182 174270 270
rect 174442 182 174830 270
rect 175002 182 175390 270
rect 175562 182 175950 270
rect 176122 182 176510 270
rect 176682 182 177070 270
rect 177242 182 177630 270
rect 177802 182 178190 270
rect 178362 182 178750 270
rect 178922 182 179310 270
rect 179482 182 179870 270
rect 180042 182 180430 270
rect 180602 182 180990 270
rect 181162 182 181550 270
rect 181722 182 182110 270
rect 182282 182 182670 270
rect 182842 182 183230 270
rect 183402 182 183790 270
rect 183962 182 184350 270
rect 184522 182 184910 270
rect 185082 182 185470 270
rect 185642 182 186030 270
rect 186202 182 186590 270
rect 186762 182 187150 270
rect 187322 182 187710 270
rect 187882 182 188270 270
rect 188442 182 188830 270
rect 189002 182 189390 270
rect 189562 182 189950 270
rect 190122 182 190510 270
rect 190682 182 191070 270
rect 191242 182 191630 270
rect 191802 182 192190 270
rect 192362 182 192750 270
rect 192922 182 193310 270
rect 193482 182 193870 270
rect 194042 182 194430 270
rect 194602 182 194990 270
rect 195162 182 195550 270
rect 195722 182 196110 270
rect 196282 182 196670 270
rect 196842 182 197230 270
rect 197402 182 197790 270
rect 197962 182 198350 270
rect 198522 182 198910 270
rect 199082 182 199470 270
rect 199642 182 200030 270
rect 200202 182 200590 270
rect 200762 182 201150 270
rect 201322 182 201710 270
rect 201882 182 202270 270
rect 202442 182 202830 270
rect 203002 182 203390 270
rect 203562 182 203950 270
rect 204122 182 204510 270
rect 204682 182 205070 270
rect 205242 182 205630 270
rect 205802 182 206190 270
rect 206362 182 206750 270
rect 206922 182 207310 270
rect 207482 182 207870 270
rect 208042 182 208430 270
rect 208602 182 208990 270
rect 209162 182 209550 270
rect 209722 182 210110 270
rect 210282 182 210670 270
rect 210842 182 211230 270
rect 211402 182 211790 270
rect 211962 182 212350 270
rect 212522 182 212910 270
rect 213082 182 213470 270
rect 213642 182 214030 270
rect 214202 182 214590 270
rect 214762 182 215150 270
rect 215322 182 215710 270
rect 215882 182 216270 270
rect 216442 182 216830 270
rect 217002 182 217390 270
rect 217562 182 217950 270
rect 218122 182 218510 270
rect 218682 182 219070 270
rect 219242 182 219630 270
rect 219802 182 220190 270
rect 220362 182 220750 270
rect 220922 182 221310 270
rect 221482 182 221870 270
rect 222042 182 222430 270
rect 222602 182 222990 270
rect 223162 182 223550 270
rect 223722 182 224110 270
rect 224282 182 224670 270
rect 224842 182 225230 270
rect 225402 182 225790 270
rect 225962 182 226350 270
rect 226522 182 226910 270
rect 227082 182 227470 270
rect 227642 182 228030 270
rect 228202 182 228590 270
rect 228762 182 229150 270
rect 229322 182 229710 270
rect 229882 182 230270 270
rect 230442 182 230830 270
rect 231002 182 231390 270
rect 231562 182 231950 270
rect 232122 182 232510 270
rect 232682 182 233070 270
rect 233242 182 233630 270
rect 233802 182 234190 270
rect 234362 182 234750 270
rect 234922 182 235310 270
rect 235482 182 235870 270
rect 236042 182 236430 270
rect 236602 182 236990 270
rect 237162 182 237550 270
rect 237722 182 238110 270
rect 238282 182 238670 270
rect 238842 182 239230 270
rect 239402 182 239790 270
rect 239962 182 240350 270
rect 240522 182 240910 270
rect 241082 182 241470 270
rect 241642 182 242030 270
rect 242202 182 242590 270
rect 242762 182 243150 270
rect 243322 182 243710 270
rect 243882 182 244270 270
rect 244442 182 244830 270
rect 245002 182 245390 270
rect 245562 182 245950 270
rect 246122 182 246510 270
rect 246682 182 247070 270
rect 247242 182 247630 270
rect 247802 182 248190 270
rect 248362 182 248750 270
rect 248922 182 249310 270
rect 249482 182 249870 270
rect 250042 182 250430 270
rect 250602 182 250990 270
rect 251162 182 251550 270
rect 251722 182 252110 270
rect 252282 182 252670 270
rect 252842 182 253230 270
rect 253402 182 253790 270
rect 253962 182 254350 270
rect 254522 182 254910 270
rect 255082 182 255470 270
rect 255642 182 256030 270
rect 256202 182 256590 270
rect 256762 182 257150 270
rect 257322 182 257710 270
rect 257882 182 258270 270
rect 258442 182 258830 270
rect 259002 182 259390 270
rect 259562 182 259950 270
rect 260122 182 260510 270
rect 260682 182 261070 270
rect 261242 182 261630 270
rect 261802 182 262190 270
rect 262362 182 262750 270
rect 262922 182 263310 270
rect 263482 182 263870 270
rect 264042 182 264430 270
rect 264602 182 264990 270
rect 265162 182 265550 270
rect 265722 182 266110 270
rect 266282 182 266670 270
rect 266842 182 267230 270
rect 267402 182 267790 270
rect 267962 182 268350 270
rect 268522 182 268910 270
rect 269082 182 269470 270
rect 269642 182 270030 270
rect 270202 182 270590 270
rect 270762 182 271150 270
rect 271322 182 271710 270
rect 271882 182 272270 270
rect 272442 182 272830 270
rect 273002 182 273390 270
rect 273562 182 273950 270
rect 274122 182 274510 270
rect 274682 182 275070 270
rect 275242 182 275630 270
rect 275802 182 276190 270
rect 276362 182 276750 270
rect 276922 182 277310 270
rect 277482 182 277870 270
rect 278042 182 278430 270
rect 278602 182 278990 270
rect 279162 182 279550 270
rect 279722 182 280110 270
rect 280282 182 280670 270
rect 280842 182 281230 270
rect 281402 182 281790 270
rect 281962 182 282350 270
rect 282522 182 282910 270
rect 283082 182 283470 270
rect 283642 182 284030 270
rect 284202 182 284590 270
rect 284762 182 285150 270
rect 285322 182 285710 270
rect 285882 182 286270 270
rect 286442 182 286830 270
rect 287002 182 287390 270
rect 287562 182 287950 270
rect 288122 182 299082 270
<< metal3 >>
rect 299760 296996 300480 297108
rect -480 296828 240 296940
rect -480 291284 240 291396
rect 299760 291340 300480 291452
rect -480 285740 240 285852
rect 299760 285684 300480 285796
rect -480 280196 240 280308
rect 299760 280028 300480 280140
rect -480 274652 240 274764
rect 299760 274372 300480 274484
rect -480 269108 240 269220
rect 299760 268716 300480 268828
rect -480 263564 240 263676
rect 299760 263060 300480 263172
rect -480 258020 240 258132
rect 299760 257404 300480 257516
rect -480 252476 240 252588
rect 299760 251748 300480 251860
rect -480 246932 240 247044
rect 299760 246092 300480 246204
rect -480 241388 240 241500
rect 299760 240436 300480 240548
rect -480 235844 240 235956
rect 299760 234780 300480 234892
rect -480 230300 240 230412
rect 299760 229124 300480 229236
rect -480 224756 240 224868
rect 299760 223468 300480 223580
rect -480 219212 240 219324
rect 299760 217812 300480 217924
rect -480 213668 240 213780
rect 299760 212156 300480 212268
rect -480 208124 240 208236
rect 299760 206500 300480 206612
rect -480 202580 240 202692
rect 299760 200844 300480 200956
rect -480 197036 240 197148
rect 299760 195188 300480 195300
rect -480 191492 240 191604
rect 299760 189532 300480 189644
rect -480 185948 240 186060
rect 299760 183876 300480 183988
rect -480 180404 240 180516
rect 299760 178220 300480 178332
rect -480 174860 240 174972
rect 299760 172564 300480 172676
rect -480 169316 240 169428
rect 299760 166908 300480 167020
rect -480 163772 240 163884
rect 299760 161252 300480 161364
rect -480 158228 240 158340
rect 299760 155596 300480 155708
rect -480 152684 240 152796
rect 299760 149940 300480 150052
rect -480 147140 240 147252
rect 299760 144284 300480 144396
rect -480 141596 240 141708
rect 299760 138628 300480 138740
rect -480 136052 240 136164
rect 299760 132972 300480 133084
rect -480 130508 240 130620
rect 299760 127316 300480 127428
rect -480 124964 240 125076
rect 299760 121660 300480 121772
rect -480 119420 240 119532
rect 299760 116004 300480 116116
rect -480 113876 240 113988
rect 299760 110348 300480 110460
rect -480 108332 240 108444
rect 299760 104692 300480 104804
rect -480 102788 240 102900
rect 299760 99036 300480 99148
rect -480 97244 240 97356
rect 299760 93380 300480 93492
rect -480 91700 240 91812
rect 299760 87724 300480 87836
rect -480 86156 240 86268
rect 299760 82068 300480 82180
rect -480 80612 240 80724
rect 299760 76412 300480 76524
rect -480 75068 240 75180
rect 299760 70756 300480 70868
rect -480 69524 240 69636
rect 299760 65100 300480 65212
rect -480 63980 240 64092
rect 299760 59444 300480 59556
rect -480 58436 240 58548
rect 299760 53788 300480 53900
rect -480 52892 240 53004
rect 299760 48132 300480 48244
rect -480 47348 240 47460
rect 299760 42476 300480 42588
rect -480 41804 240 41916
rect 299760 36820 300480 36932
rect -480 36260 240 36372
rect 299760 31164 300480 31276
rect -480 30716 240 30828
rect 299760 25508 300480 25620
rect -480 25172 240 25284
rect 299760 19852 300480 19964
rect -480 19628 240 19740
rect -480 14084 240 14196
rect 299760 14196 300480 14308
rect -480 8540 240 8652
rect 299760 8540 300480 8652
rect -480 2996 240 3108
rect 299760 2884 300480 2996
<< obsm3 >>
rect 196 297138 299810 299978
rect 196 296970 299730 297138
rect 270 296966 299730 296970
rect 270 296798 299810 296966
rect 196 291482 299810 296798
rect 196 291426 299730 291482
rect 270 291310 299730 291426
rect 270 291254 299810 291310
rect 196 285882 299810 291254
rect 270 285826 299810 285882
rect 270 285710 299730 285826
rect 196 285654 299730 285710
rect 196 280338 299810 285654
rect 270 280170 299810 280338
rect 270 280166 299730 280170
rect 196 279998 299730 280166
rect 196 274794 299810 279998
rect 270 274622 299810 274794
rect 196 274514 299810 274622
rect 196 274342 299730 274514
rect 196 269250 299810 274342
rect 270 269078 299810 269250
rect 196 268858 299810 269078
rect 196 268686 299730 268858
rect 196 263706 299810 268686
rect 270 263534 299810 263706
rect 196 263202 299810 263534
rect 196 263030 299730 263202
rect 196 258162 299810 263030
rect 270 257990 299810 258162
rect 196 257546 299810 257990
rect 196 257374 299730 257546
rect 196 252618 299810 257374
rect 270 252446 299810 252618
rect 196 251890 299810 252446
rect 196 251718 299730 251890
rect 196 247074 299810 251718
rect 270 246902 299810 247074
rect 196 246234 299810 246902
rect 196 246062 299730 246234
rect 196 241530 299810 246062
rect 270 241358 299810 241530
rect 196 240578 299810 241358
rect 196 240406 299730 240578
rect 196 235986 299810 240406
rect 270 235814 299810 235986
rect 196 234922 299810 235814
rect 196 234750 299730 234922
rect 196 230442 299810 234750
rect 270 230270 299810 230442
rect 196 229266 299810 230270
rect 196 229094 299730 229266
rect 196 224898 299810 229094
rect 270 224726 299810 224898
rect 196 223610 299810 224726
rect 196 223438 299730 223610
rect 196 219354 299810 223438
rect 270 219182 299810 219354
rect 196 217954 299810 219182
rect 196 217782 299730 217954
rect 196 213810 299810 217782
rect 270 213638 299810 213810
rect 196 212298 299810 213638
rect 196 212126 299730 212298
rect 196 208266 299810 212126
rect 270 208094 299810 208266
rect 196 206642 299810 208094
rect 196 206470 299730 206642
rect 196 202722 299810 206470
rect 270 202550 299810 202722
rect 196 200986 299810 202550
rect 196 200814 299730 200986
rect 196 197178 299810 200814
rect 270 197006 299810 197178
rect 196 195330 299810 197006
rect 196 195158 299730 195330
rect 196 191634 299810 195158
rect 270 191462 299810 191634
rect 196 189674 299810 191462
rect 196 189502 299730 189674
rect 196 186090 299810 189502
rect 270 185918 299810 186090
rect 196 184018 299810 185918
rect 196 183846 299730 184018
rect 196 180546 299810 183846
rect 270 180374 299810 180546
rect 196 178362 299810 180374
rect 196 178190 299730 178362
rect 196 175002 299810 178190
rect 270 174830 299810 175002
rect 196 172706 299810 174830
rect 196 172534 299730 172706
rect 196 169458 299810 172534
rect 270 169286 299810 169458
rect 196 167050 299810 169286
rect 196 166878 299730 167050
rect 196 163914 299810 166878
rect 270 163742 299810 163914
rect 196 161394 299810 163742
rect 196 161222 299730 161394
rect 196 158370 299810 161222
rect 270 158198 299810 158370
rect 196 155738 299810 158198
rect 196 155566 299730 155738
rect 196 152826 299810 155566
rect 270 152654 299810 152826
rect 196 150082 299810 152654
rect 196 149910 299730 150082
rect 196 147282 299810 149910
rect 270 147110 299810 147282
rect 196 144426 299810 147110
rect 196 144254 299730 144426
rect 196 141738 299810 144254
rect 270 141566 299810 141738
rect 196 138770 299810 141566
rect 196 138598 299730 138770
rect 196 136194 299810 138598
rect 270 136022 299810 136194
rect 196 133114 299810 136022
rect 196 132942 299730 133114
rect 196 130650 299810 132942
rect 270 130478 299810 130650
rect 196 127458 299810 130478
rect 196 127286 299730 127458
rect 196 125106 299810 127286
rect 270 124934 299810 125106
rect 196 121802 299810 124934
rect 196 121630 299730 121802
rect 196 119562 299810 121630
rect 270 119390 299810 119562
rect 196 116146 299810 119390
rect 196 115974 299730 116146
rect 196 114018 299810 115974
rect 270 113846 299810 114018
rect 196 110490 299810 113846
rect 196 110318 299730 110490
rect 196 108474 299810 110318
rect 270 108302 299810 108474
rect 196 104834 299810 108302
rect 196 104662 299730 104834
rect 196 102930 299810 104662
rect 270 102758 299810 102930
rect 196 99178 299810 102758
rect 196 99006 299730 99178
rect 196 97386 299810 99006
rect 270 97214 299810 97386
rect 196 93522 299810 97214
rect 196 93350 299730 93522
rect 196 91842 299810 93350
rect 270 91670 299810 91842
rect 196 87866 299810 91670
rect 196 87694 299730 87866
rect 196 86298 299810 87694
rect 270 86126 299810 86298
rect 196 82210 299810 86126
rect 196 82038 299730 82210
rect 196 80754 299810 82038
rect 270 80582 299810 80754
rect 196 76554 299810 80582
rect 196 76382 299730 76554
rect 196 75210 299810 76382
rect 270 75038 299810 75210
rect 196 70898 299810 75038
rect 196 70726 299730 70898
rect 196 69666 299810 70726
rect 270 69494 299810 69666
rect 196 65242 299810 69494
rect 196 65070 299730 65242
rect 196 64122 299810 65070
rect 270 63950 299810 64122
rect 196 59586 299810 63950
rect 196 59414 299730 59586
rect 196 58578 299810 59414
rect 270 58406 299810 58578
rect 196 53930 299810 58406
rect 196 53758 299730 53930
rect 196 53034 299810 53758
rect 270 52862 299810 53034
rect 196 48274 299810 52862
rect 196 48102 299730 48274
rect 196 47490 299810 48102
rect 270 47318 299810 47490
rect 196 42618 299810 47318
rect 196 42446 299730 42618
rect 196 41946 299810 42446
rect 270 41774 299810 41946
rect 196 36962 299810 41774
rect 196 36790 299730 36962
rect 196 36402 299810 36790
rect 270 36230 299810 36402
rect 196 31306 299810 36230
rect 196 31134 299730 31306
rect 196 30858 299810 31134
rect 270 30686 299810 30858
rect 196 25650 299810 30686
rect 196 25478 299730 25650
rect 196 25314 299810 25478
rect 270 25142 299810 25314
rect 196 19994 299810 25142
rect 196 19822 299730 19994
rect 196 19770 299810 19822
rect 270 19598 299810 19770
rect 196 14338 299810 19598
rect 196 14226 299730 14338
rect 270 14166 299730 14226
rect 270 14054 299810 14166
rect 196 8682 299810 14054
rect 270 8510 299730 8682
rect 196 3138 299810 8510
rect 270 3026 299810 3138
rect 270 2966 299730 3026
rect 196 2854 299730 2966
rect 196 854 299810 2854
<< metal4 >>
rect -11768 -10872 -11458 310752
rect -10213 -9317 -9903 309197
rect -8658 -7762 -8348 307642
rect -7103 -6207 -6793 306087
rect -5548 -4652 -5238 304532
rect -3993 -3097 -3683 302977
rect -2438 -1542 -2128 301422
rect -883 13 -573 299867
rect 2149 -10872 2459 310752
rect 4009 -10872 4319 310752
rect 5869 -10872 6179 310752
rect 7729 -10872 8039 310752
rect 9589 -10872 9899 310752
rect 11449 -10872 11759 310752
rect 13309 -10872 13619 310752
rect 15169 -10872 15479 310752
rect 17509 -10872 17819 310752
rect 19369 -10872 19679 310752
rect 21229 -10872 21539 310752
rect 23089 -10872 23399 310752
rect 24949 -10872 25259 310752
rect 26809 -10872 27119 310752
rect 28669 -10872 28979 310752
rect 30529 -10872 30839 310752
rect 32869 -10872 33179 310752
rect 34729 -10872 35039 310752
rect 36589 -10872 36899 310752
rect 38449 -10872 38759 310752
rect 40309 -10872 40619 310752
rect 42169 -10872 42479 310752
rect 44029 -10872 44339 310752
rect 45889 -10872 46199 310752
rect 48229 -10872 48539 310752
rect 50089 -10872 50399 310752
rect 51949 -10872 52259 310752
rect 53809 -10872 54119 310752
rect 55669 -10872 55979 310752
rect 57529 -10872 57839 310752
rect 59389 -10872 59699 310752
rect 61249 -10872 61559 310752
rect 63589 -10872 63899 310752
rect 65449 -10872 65759 310752
rect 67309 -10872 67619 310752
rect 69169 -10872 69479 310752
rect 71029 -10872 71339 310752
rect 72889 -10872 73199 310752
rect 74749 -10872 75059 310752
rect 76609 -10872 76919 310752
rect 78949 -10872 79259 310752
rect 80809 -10872 81119 310752
rect 82669 -10872 82979 310752
rect 84529 -10872 84839 310752
rect 86389 -10872 86699 310752
rect 88249 -10872 88559 310752
rect 90109 -10872 90419 310752
rect 91969 -10872 92279 310752
rect 94309 -10872 94619 310752
rect 96169 -10872 96479 310752
rect 98029 -10872 98339 310752
rect 99889 -10872 100199 310752
rect 101749 -10872 102059 310752
rect 103609 -10872 103919 310752
rect 105469 -10872 105779 310752
rect 107329 -10872 107639 310752
rect 109669 -10872 109979 310752
rect 111529 -10872 111839 310752
rect 113389 -10872 113699 310752
rect 115249 -10872 115559 310752
rect 117109 -10872 117419 310752
rect 118969 -10872 119279 310752
rect 120829 -10872 121139 310752
rect 122689 -10872 122999 310752
rect 125029 -10872 125339 310752
rect 126889 -10872 127199 310752
rect 128749 -10872 129059 310752
rect 130609 -10872 130919 310752
rect 132469 -10872 132779 310752
rect 134329 -10872 134639 310752
rect 136189 -10872 136499 310752
rect 138049 -10872 138359 310752
rect 140389 -10872 140699 310752
rect 142249 -10872 142559 310752
rect 144109 -10872 144419 310752
rect 145969 -10872 146279 310752
rect 147829 -10872 148139 310752
rect 149689 -10872 149999 310752
rect 151549 -10872 151859 310752
rect 153409 -10872 153719 310752
rect 155749 -10872 156059 310752
rect 157609 -10872 157919 310752
rect 159469 -10872 159779 310752
rect 161329 -10872 161639 310752
rect 163189 -10872 163499 310752
rect 165049 -10872 165359 310752
rect 166909 -10872 167219 310752
rect 168769 -10872 169079 310752
rect 171109 -10872 171419 310752
rect 172969 -10872 173279 310752
rect 174829 -10872 175139 310752
rect 176689 -10872 176999 310752
rect 178549 -10872 178859 310752
rect 180409 -10872 180719 310752
rect 182269 -10872 182579 310752
rect 184129 -10872 184439 310752
rect 186469 -10872 186779 310752
rect 188329 -10872 188639 310752
rect 190189 -10872 190499 310752
rect 192049 -10872 192359 310752
rect 193909 -10872 194219 310752
rect 195769 -10872 196079 310752
rect 197629 -10872 197939 310752
rect 199489 -10872 199799 310752
rect 201829 -10872 202139 310752
rect 203689 -10872 203999 310752
rect 205549 -10872 205859 310752
rect 207409 -10872 207719 310752
rect 209269 -10872 209579 310752
rect 211129 -10872 211439 310752
rect 212989 -10872 213299 310752
rect 214849 -10872 215159 310752
rect 217189 -10872 217499 310752
rect 219049 -10872 219359 310752
rect 220909 -10872 221219 310752
rect 222769 -10872 223079 310752
rect 224629 -10872 224939 310752
rect 226489 -10872 226799 310752
rect 228349 -10872 228659 310752
rect 230209 -10872 230519 310752
rect 232549 -10872 232859 310752
rect 234409 -10872 234719 310752
rect 236269 -10872 236579 310752
rect 238129 -10872 238439 310752
rect 239989 -10872 240299 310752
rect 241849 -10872 242159 310752
rect 243709 -10872 244019 310752
rect 245569 -10872 245879 310752
rect 247909 -10872 248219 310752
rect 249769 -10872 250079 310752
rect 251629 -10872 251939 310752
rect 253489 -10872 253799 310752
rect 255349 -10872 255659 310752
rect 257209 -10872 257519 310752
rect 259069 -10872 259379 310752
rect 260929 -10872 261239 310752
rect 263269 -10872 263579 310752
rect 265129 -10872 265439 310752
rect 266989 -10872 267299 310752
rect 268849 -10872 269159 310752
rect 270709 -10872 271019 310752
rect 272569 -10872 272879 310752
rect 274429 -10872 274739 310752
rect 276289 -10872 276599 310752
rect 278629 -10872 278939 310752
rect 280489 -10872 280799 310752
rect 282349 -10872 282659 310752
rect 284209 -10872 284519 310752
rect 286069 -10872 286379 310752
rect 287929 -10872 288239 310752
rect 289789 -10872 290099 310752
rect 291649 -10872 291959 310752
rect 293989 -10872 294299 310752
rect 295849 -10872 296159 310752
rect 297709 -10872 298019 310752
rect 300565 13 300875 299867
rect 302120 -1542 302430 301422
rect 303675 -3097 303985 302977
rect 305230 -4652 305540 304532
rect 306785 -6207 307095 306087
rect 308340 -7762 308650 307642
rect 309895 -9317 310205 309197
rect 311450 -10872 311760 310752
<< obsm4 >>
rect 14182 87481 15139 299983
rect 15509 87481 17479 299983
rect 17849 87481 19339 299983
rect 19709 87481 21199 299983
rect 21569 87481 23059 299983
rect 23429 87481 24919 299983
rect 25289 87481 26779 299983
rect 27149 87481 28639 299983
rect 29009 87481 30499 299983
rect 30869 87481 32839 299983
rect 33209 87481 34699 299983
rect 35069 87481 36559 299983
rect 36929 87481 38419 299983
rect 38789 87481 40279 299983
rect 40649 87481 42139 299983
rect 42509 87481 43999 299983
rect 44369 87481 45859 299983
rect 46229 87481 48199 299983
rect 48569 87481 50059 299983
rect 50429 87481 51919 299983
rect 52289 87481 53779 299983
rect 54149 87481 55639 299983
rect 56009 87481 57499 299983
rect 57869 87481 59359 299983
rect 59729 87481 61219 299983
rect 61589 87481 63559 299983
rect 63929 87481 65419 299983
rect 65789 87481 67279 299983
rect 67649 87481 69139 299983
rect 69509 87481 70999 299983
rect 71369 87481 72859 299983
rect 73229 87481 74719 299983
rect 75089 87481 76579 299983
rect 76949 87481 78919 299983
rect 79289 87481 80779 299983
rect 81149 87481 82639 299983
rect 83009 87481 84499 299983
rect 84869 87481 86359 299983
rect 86729 87481 88219 299983
rect 88589 87481 90079 299983
rect 90449 87481 91939 299983
rect 92309 87481 94279 299983
rect 94649 87481 96139 299983
rect 96509 87481 97999 299983
rect 98369 87481 99859 299983
rect 100229 87481 101719 299983
rect 102089 87481 103579 299983
rect 103949 87481 105439 299983
rect 105809 87481 107299 299983
rect 107669 87481 109639 299983
rect 110009 87481 111499 299983
rect 111869 87481 113359 299983
rect 113729 87481 115219 299983
rect 115589 87481 117079 299983
rect 117449 87481 118939 299983
rect 119309 87481 120799 299983
rect 121169 87481 122659 299983
rect 123029 87481 124999 299983
rect 125369 87481 126859 299983
rect 127229 87481 128719 299983
rect 129089 87481 130579 299983
rect 130949 87481 132439 299983
rect 132809 87481 134299 299983
rect 134669 87481 136159 299983
rect 136529 87481 138019 299983
rect 138389 87481 140359 299983
rect 140729 87481 142219 299983
rect 142589 87481 144079 299983
rect 144449 87481 145939 299983
rect 146309 87481 147799 299983
rect 148169 87481 149659 299983
rect 150029 87481 151519 299983
rect 151889 87481 153379 299983
rect 153749 87481 155719 299983
rect 156089 87481 157579 299983
rect 157949 87481 159439 299983
rect 159809 87481 161299 299983
rect 161669 87481 163159 299983
rect 163529 87481 165019 299983
rect 165389 87481 166879 299983
rect 167249 87481 168739 299983
rect 169109 87481 171079 299983
rect 171449 87481 172939 299983
rect 173309 87481 174799 299983
rect 175169 87481 176659 299983
rect 177029 87481 178519 299983
rect 178889 87481 180379 299983
rect 180749 87481 182239 299983
rect 182609 87481 184099 299983
rect 184469 87481 186439 299983
rect 186809 87481 188299 299983
rect 188669 87481 190159 299983
rect 190529 87481 192019 299983
rect 192389 87481 193879 299983
rect 194249 87481 195739 299983
rect 196109 87481 197599 299983
rect 197969 87481 199459 299983
rect 199829 87481 201799 299983
rect 202169 87481 203659 299983
rect 204029 87481 205519 299983
rect 205889 87481 207379 299983
rect 207749 87481 209239 299983
rect 209609 87481 211099 299983
rect 211469 87481 212959 299983
rect 213329 87481 214819 299983
rect 215189 87481 217159 299983
rect 217529 87481 219019 299983
rect 219389 87481 220879 299983
rect 221249 87481 222739 299983
rect 223109 87481 224599 299983
rect 224969 87481 226459 299983
rect 226829 87481 228319 299983
rect 228689 87481 230179 299983
rect 230549 87481 232519 299983
rect 232889 87481 234379 299983
rect 234749 87481 236239 299983
rect 236609 87481 238099 299983
rect 238469 87481 239959 299983
rect 240329 87481 241819 299983
rect 242189 87481 243679 299983
rect 244049 87481 245539 299983
rect 245909 87481 247879 299983
rect 248249 87481 249739 299983
rect 250109 87481 251599 299983
rect 251969 87481 253459 299983
rect 253829 87481 255319 299983
rect 255689 87481 257179 299983
rect 257549 87481 259039 299983
rect 259409 87481 260899 299983
rect 261269 87481 263239 299983
rect 263609 87481 265099 299983
rect 265469 87481 266959 299983
rect 267329 87481 268819 299983
rect 269189 87481 270679 299983
rect 271049 87481 272539 299983
rect 272909 87481 274399 299983
rect 274769 87481 276259 299983
rect 276629 87481 278599 299983
rect 278969 87481 280459 299983
rect 280829 87481 282319 299983
rect 282689 87481 284179 299983
rect 284549 87481 286039 299983
rect 286409 87481 287899 299983
rect 288269 87481 289759 299983
rect 290129 87481 291619 299983
rect 291989 87481 293959 299983
rect 294329 87481 295819 299983
rect 296189 87481 297679 299983
rect 298049 87481 298466 299983
<< metal5 >>
rect -11768 310442 311760 310752
rect -10213 308887 310205 309197
rect -8658 307332 308650 307642
rect -7103 305777 307095 306087
rect -5548 304222 305540 304532
rect -3993 302667 303985 302977
rect -2438 301112 302430 301422
rect -883 299557 300875 299867
rect -11768 297840 311760 298150
rect -11768 295980 311760 296290
rect -11768 294120 311760 294430
rect -11768 291822 311760 292132
rect -11768 289962 311760 290272
rect -11768 288102 311760 288412
rect -11768 286242 311760 286552
rect -11768 284382 311760 284692
rect -11768 282522 311760 282832
rect -11768 280662 311760 280972
rect -11768 278802 311760 279112
rect -11768 276504 311760 276814
rect -11768 274644 311760 274954
rect -11768 272784 311760 273094
rect -11768 270924 311760 271234
rect -11768 269064 311760 269374
rect -11768 267204 311760 267514
rect -11768 265344 311760 265654
rect -11768 263484 311760 263794
rect -11768 261186 311760 261496
rect -11768 259326 311760 259636
rect -11768 257466 311760 257776
rect -11768 255606 311760 255916
rect -11768 253746 311760 254056
rect -11768 251886 311760 252196
rect -11768 250026 311760 250336
rect -11768 248166 311760 248476
rect -11768 245868 311760 246178
rect -11768 244008 311760 244318
rect -11768 242148 311760 242458
rect -11768 240288 311760 240598
rect -11768 238428 311760 238738
rect -11768 236568 311760 236878
rect -11768 234708 311760 235018
rect -11768 232848 311760 233158
rect -11768 230550 311760 230860
rect -11768 228690 311760 229000
rect -11768 226830 311760 227140
rect -11768 224970 311760 225280
rect -11768 223110 311760 223420
rect -11768 221250 311760 221560
rect -11768 219390 311760 219700
rect -11768 217530 311760 217840
rect -11768 215232 311760 215542
rect -11768 213372 311760 213682
rect -11768 211512 311760 211822
rect -11768 209652 311760 209962
rect -11768 207792 311760 208102
rect -11768 205932 311760 206242
rect -11768 204072 311760 204382
rect -11768 202212 311760 202522
rect -11768 199914 311760 200224
rect -11768 198054 311760 198364
rect -11768 196194 311760 196504
rect -11768 194334 311760 194644
rect -11768 192474 311760 192784
rect -11768 190614 311760 190924
rect -11768 188754 311760 189064
rect -11768 186894 311760 187204
rect -11768 184596 311760 184906
rect -11768 182736 311760 183046
rect -11768 180876 311760 181186
rect -11768 179016 311760 179326
rect -11768 177156 311760 177466
rect -11768 175296 311760 175606
rect -11768 173436 311760 173746
rect -11768 171576 311760 171886
rect -11768 169278 311760 169588
rect -11768 167418 311760 167728
rect -11768 165558 311760 165868
rect -11768 163698 311760 164008
rect -11768 161838 311760 162148
rect -11768 159978 311760 160288
rect -11768 158118 311760 158428
rect -11768 156258 311760 156568
rect -11768 153960 311760 154270
rect -11768 152100 311760 152410
rect -11768 150240 311760 150550
rect -11768 148380 311760 148690
rect -11768 146520 311760 146830
rect -11768 144660 311760 144970
rect -11768 142800 311760 143110
rect -11768 140940 311760 141250
rect -11768 138642 311760 138952
rect -11768 136782 311760 137092
rect -11768 134922 311760 135232
rect -11768 133062 311760 133372
rect -11768 131202 311760 131512
rect -11768 129342 311760 129652
rect -11768 127482 311760 127792
rect -11768 125622 311760 125932
rect -11768 123324 311760 123634
rect -11768 121464 311760 121774
rect -11768 119604 311760 119914
rect -11768 117744 311760 118054
rect -11768 115884 311760 116194
rect -11768 114024 311760 114334
rect -11768 112164 311760 112474
rect -11768 110304 311760 110614
rect -11768 108006 311760 108316
rect -11768 106146 311760 106456
rect -11768 104286 311760 104596
rect -11768 102426 311760 102736
rect -11768 100566 311760 100876
rect -11768 98706 311760 99016
rect -11768 96846 311760 97156
rect -11768 94986 311760 95296
rect -11768 92688 311760 92998
rect -11768 90828 311760 91138
rect -11768 88968 311760 89278
rect -11768 87108 311760 87418
rect -11768 85248 311760 85558
rect -11768 83388 311760 83698
rect -11768 81528 311760 81838
rect -11768 79668 311760 79978
rect -11768 77370 311760 77680
rect -11768 75510 311760 75820
rect -11768 73650 311760 73960
rect -11768 71790 311760 72100
rect -11768 69930 311760 70240
rect -11768 68070 311760 68380
rect -11768 66210 311760 66520
rect -11768 64350 311760 64660
rect -11768 62052 311760 62362
rect -11768 60192 311760 60502
rect -11768 58332 311760 58642
rect -11768 56472 311760 56782
rect -11768 54612 311760 54922
rect -11768 52752 311760 53062
rect -11768 50892 311760 51202
rect -11768 49032 311760 49342
rect -11768 46734 311760 47044
rect -11768 44874 311760 45184
rect -11768 43014 311760 43324
rect -11768 41154 311760 41464
rect -11768 39294 311760 39604
rect -11768 37434 311760 37744
rect -11768 35574 311760 35884
rect -11768 33714 311760 34024
rect -11768 31416 311760 31726
rect -11768 29556 311760 29866
rect -11768 27696 311760 28006
rect -11768 25836 311760 26146
rect -11768 23976 311760 24286
rect -11768 22116 311760 22426
rect -11768 20256 311760 20566
rect -11768 18396 311760 18706
rect -11768 16098 311760 16408
rect -11768 14238 311760 14548
rect -11768 12378 311760 12688
rect -11768 10518 311760 10828
rect -11768 8658 311760 8968
rect -11768 6798 311760 7108
rect -11768 4938 311760 5248
rect -11768 3078 311760 3388
rect -883 13 300875 323
rect -2438 -1542 302430 -1232
rect -3993 -3097 303985 -2787
rect -5548 -4652 305540 -4342
rect -7103 -6207 307095 -5897
rect -8658 -7762 308650 -7452
rect -10213 -9317 310205 -9007
rect -11768 -10872 311760 -10562
<< obsm5 >>
rect 14174 298200 298474 299034
rect 14174 296340 298474 297790
rect 14174 294480 298474 295930
rect 14174 292182 298474 294070
rect 14174 290322 298474 291772
rect 14174 288462 298474 289912
rect 14174 286602 298474 288052
rect 14174 284742 298474 286192
rect 14174 282882 298474 284332
rect 14174 281022 298474 282472
rect 14174 279162 298474 280612
rect 14174 276864 298474 278752
rect 14174 275004 298474 276454
rect 14174 273144 298474 274594
rect 14174 271284 298474 272734
rect 14174 269424 298474 270874
rect 14174 267564 298474 269014
rect 14174 265704 298474 267154
rect 14174 263844 298474 265294
rect 14174 261546 298474 263434
rect 14174 259686 298474 261136
rect 14174 257826 298474 259276
rect 14174 255966 298474 257416
rect 14174 254106 298474 255556
rect 14174 252246 298474 253696
rect 14174 250386 298474 251836
rect 14174 248526 298474 249976
rect 14174 246228 298474 248116
rect 14174 244368 298474 245818
rect 14174 242508 298474 243958
rect 14174 240648 298474 242098
rect 14174 238788 298474 240238
rect 14174 236928 298474 238378
rect 14174 235068 298474 236518
rect 14174 233208 298474 234658
rect 14174 230910 298474 232798
rect 14174 229050 298474 230500
rect 14174 227190 298474 228640
rect 14174 225330 298474 226780
rect 14174 223470 298474 224920
rect 14174 221610 298474 223060
rect 14174 219750 298474 221200
rect 14174 217890 298474 219340
rect 14174 215592 298474 217480
rect 14174 213732 298474 215182
rect 14174 211872 298474 213322
rect 14174 210012 298474 211462
rect 14174 208152 298474 209602
rect 14174 206292 298474 207742
rect 14174 204432 298474 205882
rect 14174 202572 298474 204022
rect 14174 200274 298474 202162
rect 14174 198414 298474 199864
rect 14174 196554 298474 198004
rect 14174 194694 298474 196144
rect 14174 192834 298474 194284
rect 14174 190974 298474 192424
rect 14174 189114 298474 190564
rect 14174 187254 298474 188704
rect 14174 184956 298474 186844
rect 14174 183096 298474 184546
rect 14174 181236 298474 182686
rect 14174 179376 298474 180826
rect 14174 177516 298474 178966
rect 14174 175656 298474 177106
rect 14174 173796 298474 175246
rect 14174 171936 298474 173386
rect 14174 169638 298474 171526
rect 14174 167778 298474 169228
rect 14174 165918 298474 167368
rect 14174 164058 298474 165508
rect 14174 162198 298474 163648
rect 14174 160338 298474 161788
rect 14174 158478 298474 159928
rect 14174 156618 298474 158068
rect 14174 154320 298474 156208
rect 14174 152460 298474 153910
rect 14174 150600 298474 152050
rect 14174 148740 298474 150190
rect 14174 146880 298474 148330
rect 14174 145020 298474 146470
rect 14174 143160 298474 144610
rect 14174 141300 298474 142750
rect 14174 139002 298474 140890
rect 14174 137142 298474 138592
rect 14174 135282 298474 136732
rect 14174 133422 298474 134872
rect 14174 131562 298474 133012
rect 14174 129702 298474 131152
rect 14174 127842 298474 129292
rect 14174 125982 298474 127432
rect 14174 125110 298474 125572
<< labels >>
rlabel metal3 s 299760 121660 300480 121772 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 228676 299760 228788 300480 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 195524 299760 195636 300480 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 162372 299760 162484 300480 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 129220 299760 129332 300480 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 96068 299760 96180 300480 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 62916 299760 63028 300480 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 29764 299760 29876 300480 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -480 296828 240 296940 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -480 274652 240 274764 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -480 252476 240 252588 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 299760 144284 300480 144396 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -480 230300 240 230412 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -480 208124 240 208236 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -480 185948 240 186060 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -480 163772 240 163884 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -480 141596 240 141708 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -480 119420 240 119532 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -480 97244 240 97356 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -480 75068 240 75180 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -480 52892 240 53004 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 299760 166908 300480 167020 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 299760 189532 300480 189644 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 299760 212156 300480 212268 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 299760 234780 300480 234892 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 299760 257404 300480 257516 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 299760 280028 300480 280140 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 294980 299760 295092 300480 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 261828 299760 261940 300480 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 299760 2884 300480 2996 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 299760 195188 300480 195300 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 299760 217812 300480 217924 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 299760 240436 300480 240548 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 299760 263060 300480 263172 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 299760 285684 300480 285796 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 286692 299760 286804 300480 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 253540 299760 253652 300480 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 220388 299760 220500 300480 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 187236 299760 187348 300480 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 154084 299760 154196 300480 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 299760 19852 300480 19964 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 120932 299760 121044 300480 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 87780 299760 87892 300480 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 54628 299760 54740 300480 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 21476 299760 21588 300480 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -480 291284 240 291396 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -480 269108 240 269220 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -480 246932 240 247044 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -480 224756 240 224868 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -480 202580 240 202692 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -480 180404 240 180516 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 299760 36820 300480 36932 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -480 158228 240 158340 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -480 136052 240 136164 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -480 113876 240 113988 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -480 91700 240 91812 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -480 69524 240 69636 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -480 47348 240 47460 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -480 30716 240 30828 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -480 14084 240 14196 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 299760 53788 300480 53900 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 299760 70756 300480 70868 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 299760 87724 300480 87836 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 299760 104692 300480 104804 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 299760 127316 300480 127428 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 299760 149940 300480 150052 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 299760 172564 300480 172676 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 299760 14196 300480 14308 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 299760 206500 300480 206612 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 299760 229124 300480 229236 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 299760 251748 300480 251860 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 299760 274372 300480 274484 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 299760 296996 300480 297108 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 270116 299760 270228 300480 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 236964 299760 237076 300480 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 203812 299760 203924 300480 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 170660 299760 170772 300480 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 137508 299760 137620 300480 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 299760 31164 300480 31276 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 104356 299760 104468 300480 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 71204 299760 71316 300480 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 38052 299760 38164 300480 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4900 299760 5012 300480 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -480 280196 240 280308 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -480 258020 240 258132 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -480 235844 240 235956 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -480 213668 240 213780 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -480 191492 240 191604 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -480 169316 240 169428 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 299760 48132 300480 48244 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -480 147140 240 147252 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -480 124964 240 125076 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -480 102788 240 102900 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -480 80612 240 80724 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -480 58436 240 58548 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -480 36260 240 36372 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -480 19628 240 19740 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -480 2996 240 3108 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 299760 65100 300480 65212 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 299760 82068 300480 82180 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 299760 99036 300480 99148 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 299760 116004 300480 116116 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 299760 138628 300480 138740 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 299760 161252 300480 161364 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 299760 183876 300480 183988 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 299760 8540 300480 8652 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 299760 200844 300480 200956 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 299760 223468 300480 223580 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 299760 246092 300480 246204 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 299760 268716 300480 268828 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 299760 291340 300480 291452 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 278404 299760 278516 300480 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 245252 299760 245364 300480 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 212100 299760 212212 300480 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 178948 299760 179060 300480 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 145796 299760 145908 300480 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 299760 25508 300480 25620 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 112644 299760 112756 300480 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 79492 299760 79604 300480 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 46340 299760 46452 300480 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 13188 299760 13300 300480 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -480 285740 240 285852 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -480 263564 240 263676 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -480 241388 240 241500 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -480 219212 240 219324 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -480 197036 240 197148 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -480 174860 240 174972 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 299760 42476 300480 42588 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -480 152684 240 152796 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -480 130508 240 130620 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -480 108332 240 108444 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -480 86156 240 86268 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -480 63980 240 64092 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -480 41804 240 41916 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -480 25172 240 25284 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -480 8540 240 8652 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 299760 59444 300480 59556 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 299760 76412 300480 76524 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 299760 93380 300480 93492 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 299760 110348 300480 110460 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 299760 132972 300480 133084 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 299760 155596 300480 155708 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 299760 178220 300480 178332 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 71260 -480 71372 240 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 239260 -480 239372 240 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 240940 -480 241052 240 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 242620 -480 242732 240 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 244300 -480 244412 240 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 245980 -480 246092 240 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 247660 -480 247772 240 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 249340 -480 249452 240 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 251020 -480 251132 240 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 252700 -480 252812 240 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 254380 -480 254492 240 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 88060 -480 88172 240 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 256060 -480 256172 240 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 257740 -480 257852 240 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 259420 -480 259532 240 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 261100 -480 261212 240 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 262780 -480 262892 240 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 264460 -480 264572 240 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 266140 -480 266252 240 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 267820 -480 267932 240 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 269500 -480 269612 240 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 271180 -480 271292 240 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 89740 -480 89852 240 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 272860 -480 272972 240 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 274540 -480 274652 240 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 276220 -480 276332 240 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 277900 -480 278012 240 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 279580 -480 279692 240 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 281260 -480 281372 240 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 282940 -480 283052 240 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 284620 -480 284732 240 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 91420 -480 91532 240 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 93100 -480 93212 240 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 94780 -480 94892 240 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 96460 -480 96572 240 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 98140 -480 98252 240 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 99820 -480 99932 240 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 101500 -480 101612 240 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 103180 -480 103292 240 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 72940 -480 73052 240 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 104860 -480 104972 240 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 106540 -480 106652 240 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 108220 -480 108332 240 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 109900 -480 110012 240 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 111580 -480 111692 240 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 113260 -480 113372 240 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 114940 -480 115052 240 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 116620 -480 116732 240 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 118300 -480 118412 240 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 119980 -480 120092 240 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 74620 -480 74732 240 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 121660 -480 121772 240 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 123340 -480 123452 240 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 125020 -480 125132 240 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 126700 -480 126812 240 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 128380 -480 128492 240 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 130060 -480 130172 240 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 131740 -480 131852 240 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 133420 -480 133532 240 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 135100 -480 135212 240 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 136780 -480 136892 240 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 76300 -480 76412 240 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 138460 -480 138572 240 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 140140 -480 140252 240 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 141820 -480 141932 240 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 143500 -480 143612 240 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 145180 -480 145292 240 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 146860 -480 146972 240 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 148540 -480 148652 240 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 150220 -480 150332 240 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 151900 -480 152012 240 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 153580 -480 153692 240 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 77980 -480 78092 240 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 155260 -480 155372 240 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 156940 -480 157052 240 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 158620 -480 158732 240 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 160300 -480 160412 240 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 161980 -480 162092 240 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 163660 -480 163772 240 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 165340 -480 165452 240 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 167020 -480 167132 240 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 168700 -480 168812 240 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 170380 -480 170492 240 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 79660 -480 79772 240 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 172060 -480 172172 240 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 173740 -480 173852 240 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 175420 -480 175532 240 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 177100 -480 177212 240 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 178780 -480 178892 240 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 180460 -480 180572 240 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 182140 -480 182252 240 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 183820 -480 183932 240 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 185500 -480 185612 240 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 187180 -480 187292 240 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 81340 -480 81452 240 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 188860 -480 188972 240 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 190540 -480 190652 240 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 192220 -480 192332 240 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 193900 -480 194012 240 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 195580 -480 195692 240 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 197260 -480 197372 240 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 198940 -480 199052 240 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 200620 -480 200732 240 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 202300 -480 202412 240 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 203980 -480 204092 240 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 83020 -480 83132 240 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 205660 -480 205772 240 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 207340 -480 207452 240 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 209020 -480 209132 240 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 210700 -480 210812 240 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 212380 -480 212492 240 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 214060 -480 214172 240 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 215740 -480 215852 240 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 217420 -480 217532 240 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 219100 -480 219212 240 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 220780 -480 220892 240 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 84700 -480 84812 240 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 222460 -480 222572 240 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 224140 -480 224252 240 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 225820 -480 225932 240 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 227500 -480 227612 240 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 229180 -480 229292 240 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 230860 -480 230972 240 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 232540 -480 232652 240 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 234220 -480 234332 240 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 235900 -480 236012 240 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 237580 -480 237692 240 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 86380 -480 86492 240 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 71820 -480 71932 240 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 239820 -480 239932 240 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 241500 -480 241612 240 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 243180 -480 243292 240 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 244860 -480 244972 240 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 246540 -480 246652 240 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 248220 -480 248332 240 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 249900 -480 250012 240 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 251580 -480 251692 240 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 253260 -480 253372 240 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 254940 -480 255052 240 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 88620 -480 88732 240 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 256620 -480 256732 240 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 258300 -480 258412 240 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 259980 -480 260092 240 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 261660 -480 261772 240 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 263340 -480 263452 240 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 265020 -480 265132 240 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 266700 -480 266812 240 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 268380 -480 268492 240 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 270060 -480 270172 240 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 271740 -480 271852 240 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 90300 -480 90412 240 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 273420 -480 273532 240 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 275100 -480 275212 240 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 276780 -480 276892 240 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 278460 -480 278572 240 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 280140 -480 280252 240 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 281820 -480 281932 240 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 283500 -480 283612 240 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 285180 -480 285292 240 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 91980 -480 92092 240 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 93660 -480 93772 240 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 95340 -480 95452 240 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 97020 -480 97132 240 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 98700 -480 98812 240 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 100380 -480 100492 240 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 102060 -480 102172 240 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 103740 -480 103852 240 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 73500 -480 73612 240 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 105420 -480 105532 240 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 107100 -480 107212 240 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 108780 -480 108892 240 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 110460 -480 110572 240 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 112140 -480 112252 240 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 113820 -480 113932 240 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 115500 -480 115612 240 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 117180 -480 117292 240 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 118860 -480 118972 240 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 120540 -480 120652 240 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 75180 -480 75292 240 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 122220 -480 122332 240 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 123900 -480 124012 240 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 125580 -480 125692 240 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 127260 -480 127372 240 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 128940 -480 129052 240 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 130620 -480 130732 240 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 132300 -480 132412 240 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 133980 -480 134092 240 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 135660 -480 135772 240 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 137340 -480 137452 240 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 76860 -480 76972 240 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 139020 -480 139132 240 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 140700 -480 140812 240 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 142380 -480 142492 240 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 144060 -480 144172 240 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 145740 -480 145852 240 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 147420 -480 147532 240 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 149100 -480 149212 240 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 150780 -480 150892 240 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 152460 -480 152572 240 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 154140 -480 154252 240 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 78540 -480 78652 240 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 155820 -480 155932 240 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 157500 -480 157612 240 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 159180 -480 159292 240 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 160860 -480 160972 240 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 162540 -480 162652 240 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 164220 -480 164332 240 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 165900 -480 166012 240 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 167580 -480 167692 240 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 169260 -480 169372 240 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 170940 -480 171052 240 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 80220 -480 80332 240 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 172620 -480 172732 240 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 174300 -480 174412 240 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 175980 -480 176092 240 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 177660 -480 177772 240 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 179340 -480 179452 240 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 181020 -480 181132 240 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 182700 -480 182812 240 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 184380 -480 184492 240 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 186060 -480 186172 240 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 187740 -480 187852 240 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 81900 -480 82012 240 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 189420 -480 189532 240 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 191100 -480 191212 240 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 192780 -480 192892 240 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 194460 -480 194572 240 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 196140 -480 196252 240 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 197820 -480 197932 240 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 199500 -480 199612 240 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 201180 -480 201292 240 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 202860 -480 202972 240 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 204540 -480 204652 240 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 83580 -480 83692 240 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 206220 -480 206332 240 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 207900 -480 208012 240 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 209580 -480 209692 240 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 211260 -480 211372 240 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 212940 -480 213052 240 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 214620 -480 214732 240 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 216300 -480 216412 240 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 217980 -480 218092 240 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 219660 -480 219772 240 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 221340 -480 221452 240 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 85260 -480 85372 240 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 223020 -480 223132 240 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 224700 -480 224812 240 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 226380 -480 226492 240 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 228060 -480 228172 240 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 229740 -480 229852 240 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 231420 -480 231532 240 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 233100 -480 233212 240 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 234780 -480 234892 240 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 236460 -480 236572 240 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 238140 -480 238252 240 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 86940 -480 87052 240 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 72380 -480 72492 240 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 240380 -480 240492 240 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 242060 -480 242172 240 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 243740 -480 243852 240 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 245420 -480 245532 240 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 247100 -480 247212 240 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 248780 -480 248892 240 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 250460 -480 250572 240 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 252140 -480 252252 240 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 253820 -480 253932 240 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 255500 -480 255612 240 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 89180 -480 89292 240 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 257180 -480 257292 240 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 258860 -480 258972 240 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 260540 -480 260652 240 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 262220 -480 262332 240 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 263900 -480 264012 240 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 265580 -480 265692 240 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 267260 -480 267372 240 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 268940 -480 269052 240 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 270620 -480 270732 240 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 272300 -480 272412 240 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 90860 -480 90972 240 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 273980 -480 274092 240 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 275660 -480 275772 240 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 277340 -480 277452 240 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 279020 -480 279132 240 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 280700 -480 280812 240 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 282380 -480 282492 240 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 284060 -480 284172 240 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 285740 -480 285852 240 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 92540 -480 92652 240 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 94220 -480 94332 240 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 95900 -480 96012 240 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 97580 -480 97692 240 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 99260 -480 99372 240 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 100940 -480 101052 240 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 102620 -480 102732 240 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 104300 -480 104412 240 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 74060 -480 74172 240 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 105980 -480 106092 240 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 107660 -480 107772 240 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 109340 -480 109452 240 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 111020 -480 111132 240 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 112700 -480 112812 240 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 114380 -480 114492 240 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 116060 -480 116172 240 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 117740 -480 117852 240 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 119420 -480 119532 240 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 121100 -480 121212 240 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 75740 -480 75852 240 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 122780 -480 122892 240 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 124460 -480 124572 240 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 126140 -480 126252 240 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 127820 -480 127932 240 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 129500 -480 129612 240 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 131180 -480 131292 240 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 132860 -480 132972 240 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 134540 -480 134652 240 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 136220 -480 136332 240 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 137900 -480 138012 240 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 77420 -480 77532 240 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 139580 -480 139692 240 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 141260 -480 141372 240 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 142940 -480 143052 240 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 144620 -480 144732 240 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 146300 -480 146412 240 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 147980 -480 148092 240 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 149660 -480 149772 240 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 151340 -480 151452 240 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 153020 -480 153132 240 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 154700 -480 154812 240 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 79100 -480 79212 240 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 156380 -480 156492 240 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 158060 -480 158172 240 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 159740 -480 159852 240 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 161420 -480 161532 240 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 163100 -480 163212 240 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 164780 -480 164892 240 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 166460 -480 166572 240 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 168140 -480 168252 240 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 169820 -480 169932 240 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 171500 -480 171612 240 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 80780 -480 80892 240 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 173180 -480 173292 240 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 174860 -480 174972 240 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 176540 -480 176652 240 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 178220 -480 178332 240 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 179900 -480 180012 240 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 181580 -480 181692 240 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 183260 -480 183372 240 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 184940 -480 185052 240 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 186620 -480 186732 240 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 188300 -480 188412 240 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 82460 -480 82572 240 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 189980 -480 190092 240 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 191660 -480 191772 240 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 193340 -480 193452 240 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 195020 -480 195132 240 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 196700 -480 196812 240 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 198380 -480 198492 240 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 200060 -480 200172 240 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 201740 -480 201852 240 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 203420 -480 203532 240 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 205100 -480 205212 240 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 84140 -480 84252 240 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 206780 -480 206892 240 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 208460 -480 208572 240 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 210140 -480 210252 240 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 211820 -480 211932 240 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 213500 -480 213612 240 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 215180 -480 215292 240 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 216860 -480 216972 240 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 218540 -480 218652 240 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 220220 -480 220332 240 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 221900 -480 222012 240 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 85820 -480 85932 240 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 223580 -480 223692 240 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 225260 -480 225372 240 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 226940 -480 227052 240 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 228620 -480 228732 240 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 230300 -480 230412 240 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 231980 -480 232092 240 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 233660 -480 233772 240 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 235340 -480 235452 240 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 237020 -480 237132 240 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 238700 -480 238812 240 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 87500 -480 87612 240 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 286300 -480 286412 240 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 286860 -480 286972 240 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 287420 -480 287532 240 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 287980 -480 288092 240 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -883 13 -573 299867 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -883 13 300875 323 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -883 299557 300875 299867 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 300565 13 300875 299867 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 2149 -10872 2459 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 17509 -10872 17819 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 32869 -10872 33179 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 48229 -10872 48539 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 63589 -10872 63899 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 78949 -10872 79259 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 94309 -10872 94619 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109669 -10872 109979 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 125029 -10872 125339 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 140389 -10872 140699 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 155749 -10872 156059 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 171109 -10872 171419 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 186469 -10872 186779 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 201829 -10872 202139 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217189 -10872 217499 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 232549 -10872 232859 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 247909 -10872 248219 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 263269 -10872 263579 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 278629 -10872 278939 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 293989 -10872 294299 310752 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 3078 311760 3388 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 18396 311760 18706 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 33714 311760 34024 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 49032 311760 49342 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 64350 311760 64660 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 79668 311760 79978 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 94986 311760 95296 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 110304 311760 110614 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 125622 311760 125932 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 140940 311760 141250 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 156258 311760 156568 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 171576 311760 171886 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 186894 311760 187204 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 202212 311760 202522 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 217530 311760 217840 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 232848 311760 233158 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 248166 311760 248476 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 263484 311760 263794 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 278802 311760 279112 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -11768 294120 311760 294430 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3993 -3097 -3683 302977 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3993 -3097 303985 -2787 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3993 302667 303985 302977 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 303675 -3097 303985 302977 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 5869 -10872 6179 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 21229 -10872 21539 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 36589 -10872 36899 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 51949 -10872 52259 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 67309 -10872 67619 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 82669 -10872 82979 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 98029 -10872 98339 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 113389 -10872 113699 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 128749 -10872 129059 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 144109 -10872 144419 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 159469 -10872 159779 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 174829 -10872 175139 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 190189 -10872 190499 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 205549 -10872 205859 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 220909 -10872 221219 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 236269 -10872 236579 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 251629 -10872 251939 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 266989 -10872 267299 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 282349 -10872 282659 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 297709 -10872 298019 310752 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 6798 311760 7108 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 22116 311760 22426 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 37434 311760 37744 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 52752 311760 53062 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 68070 311760 68380 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 83388 311760 83698 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 98706 311760 99016 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 114024 311760 114334 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 129342 311760 129652 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 144660 311760 144970 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 159978 311760 160288 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 175296 311760 175606 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 190614 311760 190924 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 205932 311760 206242 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 221250 311760 221560 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 236568 311760 236878 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 251886 311760 252196 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 267204 311760 267514 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 282522 311760 282832 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -11768 297840 311760 298150 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -7103 -6207 -6793 306087 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -7103 -6207 307095 -5897 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -7103 305777 307095 306087 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 306785 -6207 307095 306087 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 9589 -10872 9899 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 24949 -10872 25259 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 40309 -10872 40619 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 55669 -10872 55979 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 71029 -10872 71339 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 86389 -10872 86699 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 101749 -10872 102059 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 117109 -10872 117419 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 132469 -10872 132779 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 147829 -10872 148139 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 163189 -10872 163499 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 178549 -10872 178859 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 193909 -10872 194219 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 209269 -10872 209579 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 224629 -10872 224939 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 239989 -10872 240299 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 255349 -10872 255659 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 270709 -10872 271019 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 286069 -10872 286379 310752 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 10518 311760 10828 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 25836 311760 26146 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 41154 311760 41464 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 56472 311760 56782 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 71790 311760 72100 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 87108 311760 87418 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 102426 311760 102736 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 117744 311760 118054 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 133062 311760 133372 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 148380 311760 148690 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 163698 311760 164008 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 179016 311760 179326 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 194334 311760 194644 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 209652 311760 209962 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 224970 311760 225280 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 240288 311760 240598 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 255606 311760 255916 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 270924 311760 271234 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -11768 286242 311760 286552 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -10213 -9317 -9903 309197 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -10213 -9317 310205 -9007 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -10213 308887 310205 309197 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 309895 -9317 310205 309197 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 13309 -10872 13619 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 28669 -10872 28979 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 44029 -10872 44339 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 59389 -10872 59699 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 74749 -10872 75059 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 90109 -10872 90419 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 105469 -10872 105779 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 120829 -10872 121139 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 136189 -10872 136499 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 151549 -10872 151859 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 166909 -10872 167219 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 182269 -10872 182579 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 197629 -10872 197939 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 212989 -10872 213299 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 228349 -10872 228659 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 243709 -10872 244019 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 259069 -10872 259379 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 274429 -10872 274739 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 289789 -10872 290099 310752 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 14238 311760 14548 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 29556 311760 29866 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 44874 311760 45184 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 60192 311760 60502 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 75510 311760 75820 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 90828 311760 91138 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 106146 311760 106456 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 121464 311760 121774 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 136782 311760 137092 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 152100 311760 152410 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 167418 311760 167728 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 182736 311760 183046 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 198054 311760 198364 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 213372 311760 213682 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 228690 311760 229000 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 244008 311760 244318 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 259326 311760 259636 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 274644 311760 274954 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -11768 289962 311760 290272 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -8658 -7762 -8348 307642 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8658 -7762 308650 -7452 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8658 307332 308650 307642 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 308340 -7762 308650 307642 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 11449 -10872 11759 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 26809 -10872 27119 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 42169 -10872 42479 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 57529 -10872 57839 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 72889 -10872 73199 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 88249 -10872 88559 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 103609 -10872 103919 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 118969 -10872 119279 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 134329 -10872 134639 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 149689 -10872 149999 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 165049 -10872 165359 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 180409 -10872 180719 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 195769 -10872 196079 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 211129 -10872 211439 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 226489 -10872 226799 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 241849 -10872 242159 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 257209 -10872 257519 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 272569 -10872 272879 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 287929 -10872 288239 310752 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 12378 311760 12688 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 27696 311760 28006 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 43014 311760 43324 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 58332 311760 58642 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 73650 311760 73960 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 88968 311760 89278 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 104286 311760 104596 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 119604 311760 119914 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 134922 311760 135232 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 150240 311760 150550 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 165558 311760 165868 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 180876 311760 181186 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 196194 311760 196504 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 211512 311760 211822 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 226830 311760 227140 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 242148 311760 242458 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 257466 311760 257776 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 272784 311760 273094 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -11768 288102 311760 288412 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -11768 -10872 -11458 310752 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 -10872 311760 -10562 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 310442 311760 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 311450 -10872 311760 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 15169 -10872 15479 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 30529 -10872 30839 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 45889 -10872 46199 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 61249 -10872 61559 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 76609 -10872 76919 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 91969 -10872 92279 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 107329 -10872 107639 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 122689 -10872 122999 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 138049 -10872 138359 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 153409 -10872 153719 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 168769 -10872 169079 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 184129 -10872 184439 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 199489 -10872 199799 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 214849 -10872 215159 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 230209 -10872 230519 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 245569 -10872 245879 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 260929 -10872 261239 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 276289 -10872 276599 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 291649 -10872 291959 310752 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 16098 311760 16408 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 31416 311760 31726 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 46734 311760 47044 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 62052 311760 62362 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 77370 311760 77680 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 92688 311760 92998 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 108006 311760 108316 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 123324 311760 123634 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 138642 311760 138952 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 153960 311760 154270 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 169278 311760 169588 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 184596 311760 184906 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 199914 311760 200224 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 215232 311760 215542 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 230550 311760 230860 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 245868 311760 246178 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 261186 311760 261496 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 276504 311760 276814 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -11768 291822 311760 292132 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2438 -1542 -2128 301422 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2438 -1542 302430 -1232 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2438 301112 302430 301422 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 302120 -1542 302430 301422 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 4009 -10872 4319 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 19369 -10872 19679 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 34729 -10872 35039 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 50089 -10872 50399 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 65449 -10872 65759 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 80809 -10872 81119 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 96169 -10872 96479 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 111529 -10872 111839 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 126889 -10872 127199 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 142249 -10872 142559 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 157609 -10872 157919 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 172969 -10872 173279 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 188329 -10872 188639 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 203689 -10872 203999 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 219049 -10872 219359 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 234409 -10872 234719 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 249769 -10872 250079 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 265129 -10872 265439 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 280489 -10872 280799 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 295849 -10872 296159 310752 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 4938 311760 5248 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 20256 311760 20566 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 35574 311760 35884 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 50892 311760 51202 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 66210 311760 66520 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 81528 311760 81838 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 96846 311760 97156 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 112164 311760 112474 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 127482 311760 127792 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 142800 311760 143110 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 158118 311760 158428 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 173436 311760 173746 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 188754 311760 189064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 204072 311760 204382 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 219390 311760 219700 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 234708 311760 235018 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 250026 311760 250336 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 265344 311760 265654 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 280662 311760 280972 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -11768 295980 311760 296290 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -5548 -4652 -5238 304532 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5548 -4652 305540 -4342 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -5548 304222 305540 304532 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 305230 -4652 305540 304532 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 7729 -10872 8039 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 23089 -10872 23399 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 38449 -10872 38759 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 53809 -10872 54119 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 69169 -10872 69479 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84529 -10872 84839 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 99889 -10872 100199 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 115249 -10872 115559 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 130609 -10872 130919 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 145969 -10872 146279 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 161329 -10872 161639 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 176689 -10872 176999 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192049 -10872 192359 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 207409 -10872 207719 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 222769 -10872 223079 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 238129 -10872 238439 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 253489 -10872 253799 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 268849 -10872 269159 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 284209 -10872 284519 310752 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 8658 311760 8968 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 23976 311760 24286 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 39294 311760 39604 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 54612 311760 54922 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 69930 311760 70240 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 85248 311760 85558 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 100566 311760 100876 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 115884 311760 116194 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 131202 311760 131512 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 146520 311760 146830 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 161838 311760 162148 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 177156 311760 177466 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 192474 311760 192784 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 207792 311760 208102 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 223110 311760 223420 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 238428 311760 238738 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 253746 311760 254056 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 269064 311760 269374 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -11768 284382 311760 284692 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 11900 -480 12012 240 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 12460 -480 12572 240 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 13020 -480 13132 240 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 15260 -480 15372 240 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 34300 -480 34412 240 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 35980 -480 36092 240 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 37660 -480 37772 240 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 39340 -480 39452 240 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 41020 -480 41132 240 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 42700 -480 42812 240 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 44380 -480 44492 240 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 46060 -480 46172 240 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 47740 -480 47852 240 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 49420 -480 49532 240 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 17500 -480 17612 240 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 51100 -480 51212 240 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 52780 -480 52892 240 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 54460 -480 54572 240 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 56140 -480 56252 240 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 57820 -480 57932 240 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 59500 -480 59612 240 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 61180 -480 61292 240 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 62860 -480 62972 240 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 64540 -480 64652 240 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 66220 -480 66332 240 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 19740 -480 19852 240 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 67900 -480 68012 240 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 69580 -480 69692 240 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21980 -480 22092 240 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 24220 -480 24332 240 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 25900 -480 26012 240 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 27580 -480 27692 240 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 29260 -480 29372 240 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 30940 -480 31052 240 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 32620 -480 32732 240 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 13580 -480 13692 240 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 15820 -480 15932 240 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 34860 -480 34972 240 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 36540 -480 36652 240 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 38220 -480 38332 240 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 39900 -480 40012 240 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 41580 -480 41692 240 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 43260 -480 43372 240 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 44940 -480 45052 240 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 46620 -480 46732 240 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 48300 -480 48412 240 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 49980 -480 50092 240 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 18060 -480 18172 240 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 51660 -480 51772 240 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 53340 -480 53452 240 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 55020 -480 55132 240 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 56700 -480 56812 240 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 58380 -480 58492 240 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 60060 -480 60172 240 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 61740 -480 61852 240 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 63420 -480 63532 240 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 65100 -480 65212 240 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 66780 -480 66892 240 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 20300 -480 20412 240 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 68460 -480 68572 240 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 70140 -480 70252 240 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22540 -480 22652 240 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 24780 -480 24892 240 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 26460 -480 26572 240 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 28140 -480 28252 240 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 29820 -480 29932 240 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 31500 -480 31612 240 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 33180 -480 33292 240 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 16380 -480 16492 240 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 35420 -480 35532 240 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 37100 -480 37212 240 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 38780 -480 38892 240 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 40460 -480 40572 240 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 42140 -480 42252 240 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 43820 -480 43932 240 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 45500 -480 45612 240 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 47180 -480 47292 240 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 48860 -480 48972 240 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 50540 -480 50652 240 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 18620 -480 18732 240 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 52220 -480 52332 240 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 53900 -480 54012 240 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 55580 -480 55692 240 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 57260 -480 57372 240 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 58940 -480 59052 240 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 60620 -480 60732 240 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 62300 -480 62412 240 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 63980 -480 64092 240 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 65660 -480 65772 240 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 67340 -480 67452 240 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 20860 -480 20972 240 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 69020 -480 69132 240 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 70700 -480 70812 240 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 23100 -480 23212 240 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 25340 -480 25452 240 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 27020 -480 27132 240 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 28700 -480 28812 240 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 30380 -480 30492 240 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 32060 -480 32172 240 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 33740 -480 33852 240 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 16940 -480 17052 240 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 19180 -480 19292 240 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 21420 -480 21532 240 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 23660 -480 23772 240 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 14140 -480 14252 240 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 14700 -480 14812 240 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 300000 300000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 133890904
string GDS_FILE /Volumes/Efabless/ParaRAM/openlane/user_project_wrapper/runs/22_11_07_11_52/results/signoff/user_project_wrapper.magic.gds
string GDS_START 320528
<< end >>

