magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -183 117 183 136
rect -183 -117 -164 117
rect 164 -117 183 117
rect -183 -136 183 -117
<< psubdiffcont >>
rect -164 -117 164 117
<< metal1 >>
rect -175 117 175 128
rect -175 -117 -164 117
rect 164 -117 175 117
rect -175 -128 175 -117
<< properties >>
string GDS_END 537116
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 536152
<< end >>
