magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -64 1876 65 1917
rect -64 1824 -26 1876
rect 26 1824 65 1876
rect -64 1658 65 1824
rect -64 1606 -26 1658
rect 26 1606 65 1658
rect -64 1441 65 1606
rect -64 1389 -26 1441
rect 26 1389 65 1441
rect -64 1223 65 1389
rect -64 1171 -26 1223
rect 26 1171 65 1223
rect -64 1005 65 1171
rect -64 953 -26 1005
rect 26 953 65 1005
rect -64 788 65 953
rect -64 736 -26 788
rect 26 736 65 788
rect -64 570 65 736
rect -64 518 -26 570
rect 26 518 65 570
rect -64 353 65 518
rect -64 301 -26 353
rect 26 301 65 353
rect -64 135 65 301
rect -64 83 -26 135
rect 26 83 65 135
rect -64 -83 65 83
rect -64 -135 -26 -83
rect 26 -135 65 -83
rect -64 -301 65 -135
rect -64 -353 -26 -301
rect 26 -353 65 -301
rect -64 -518 65 -353
rect -64 -570 -26 -518
rect 26 -570 65 -518
rect -64 -736 65 -570
rect -64 -788 -26 -736
rect 26 -788 65 -736
rect -64 -953 65 -788
rect -64 -1005 -26 -953
rect 26 -1005 65 -953
rect -64 -1171 65 -1005
rect -64 -1223 -26 -1171
rect 26 -1223 65 -1171
rect -64 -1389 65 -1223
rect -64 -1441 -26 -1389
rect 26 -1441 65 -1389
rect -64 -1606 65 -1441
rect -64 -1658 -26 -1606
rect 26 -1658 65 -1606
rect -64 -1824 65 -1658
rect -64 -1876 -26 -1824
rect 26 -1876 65 -1824
rect -64 -1916 65 -1876
rect -57 -1917 58 -1916
<< via1 >>
rect -26 1824 26 1876
rect -26 1606 26 1658
rect -26 1389 26 1441
rect -26 1171 26 1223
rect -26 953 26 1005
rect -26 736 26 788
rect -26 518 26 570
rect -26 301 26 353
rect -26 83 26 135
rect -26 -135 26 -83
rect -26 -353 26 -301
rect -26 -570 26 -518
rect -26 -788 26 -736
rect -26 -1005 26 -953
rect -26 -1223 26 -1171
rect -26 -1441 26 -1389
rect -26 -1658 26 -1606
rect -26 -1876 26 -1824
<< metal2 >>
rect -64 1876 65 1917
rect -64 1824 -26 1876
rect 26 1824 65 1876
rect -64 1658 65 1824
rect -64 1606 -26 1658
rect 26 1606 65 1658
rect -64 1441 65 1606
rect -64 1389 -26 1441
rect 26 1389 65 1441
rect -64 1223 65 1389
rect -64 1171 -26 1223
rect 26 1171 65 1223
rect -64 1005 65 1171
rect -64 953 -26 1005
rect 26 953 65 1005
rect -64 788 65 953
rect -64 736 -26 788
rect 26 736 65 788
rect -64 570 65 736
rect -64 518 -26 570
rect 26 518 65 570
rect -64 353 65 518
rect -64 301 -26 353
rect 26 301 65 353
rect -64 135 65 301
rect -64 83 -26 135
rect 26 83 65 135
rect -64 -83 65 83
rect -64 -135 -26 -83
rect 26 -135 65 -83
rect -64 -301 65 -135
rect -64 -353 -26 -301
rect 26 -353 65 -301
rect -64 -518 65 -353
rect -64 -570 -26 -518
rect 26 -570 65 -518
rect -64 -736 65 -570
rect -64 -788 -26 -736
rect 26 -788 65 -736
rect -64 -953 65 -788
rect -64 -1005 -26 -953
rect 26 -1005 65 -953
rect -64 -1171 65 -1005
rect -64 -1223 -26 -1171
rect 26 -1223 65 -1171
rect -64 -1389 65 -1223
rect -64 -1441 -26 -1389
rect 26 -1441 65 -1389
rect -64 -1606 65 -1441
rect -64 -1658 -26 -1606
rect 26 -1658 65 -1606
rect -64 -1824 65 -1658
rect -64 -1876 -26 -1824
rect 26 -1876 65 -1824
rect -64 -1916 65 -1876
<< properties >>
string GDS_END 1037678
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1036362
<< end >>
