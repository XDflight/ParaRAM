magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 44323 242 44342
rect -42 -23 -23 44323
rect 223 -23 242 44323
rect -42 -42 242 -23
<< psubdiffcont >>
rect -23 -23 223 44323
<< metal1 >>
rect -34 44323 234 44334
rect -34 -23 -23 44323
rect 223 -23 234 44323
rect -34 -34 234 -23
<< properties >>
string GDS_END 1733242
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1647798
<< end >>
