magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 4902 1094
<< pwell >>
rect -86 -86 4902 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 732 215 852 333
rect 956 215 1076 333
rect 1180 215 1300 333
rect 1348 215 1468 333
rect 1580 215 1700 333
rect 1804 215 1924 333
rect 1972 215 2092 333
rect 2196 215 2316 333
rect 2420 215 2540 333
rect 2964 175 3084 333
rect 3132 175 3252 333
rect 3356 175 3476 333
rect 3524 175 3644 333
rect 3892 69 4012 333
rect 4116 69 4236 333
rect 4340 69 4460 333
rect 4564 69 4684 333
<< mvpmos >>
rect 124 573 224 849
rect 328 573 428 849
rect 676 573 776 773
rect 880 573 980 773
rect 1084 573 1184 773
rect 1288 573 1388 773
rect 1580 690 1680 890
rect 1928 690 2028 890
rect 2208 573 2308 773
rect 2412 573 2512 773
rect 2616 573 2716 773
rect 2964 573 3064 849
rect 3168 573 3268 849
rect 3372 573 3472 849
rect 3576 573 3676 849
rect 3924 573 4024 939
rect 4128 573 4228 939
rect 4332 573 4432 939
rect 4536 573 4636 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 468 175 556 274
rect 644 274 732 333
rect 644 228 657 274
rect 703 228 732 274
rect 644 215 732 228
rect 852 320 956 333
rect 852 274 881 320
rect 927 274 956 320
rect 852 215 956 274
rect 1076 320 1180 333
rect 1076 274 1105 320
rect 1151 274 1180 320
rect 1076 215 1180 274
rect 1300 215 1348 333
rect 1468 215 1580 333
rect 1700 274 1804 333
rect 1700 228 1729 274
rect 1775 228 1804 274
rect 1700 215 1804 228
rect 1924 215 1972 333
rect 2092 320 2196 333
rect 2092 274 2121 320
rect 2167 274 2196 320
rect 2092 215 2196 274
rect 2316 320 2420 333
rect 2316 274 2345 320
rect 2391 274 2420 320
rect 2316 215 2420 274
rect 2540 319 2628 333
rect 2540 273 2569 319
rect 2615 273 2628 319
rect 2540 215 2628 273
rect 2876 297 2964 333
rect 2876 251 2889 297
rect 2935 251 2964 297
rect 2876 175 2964 251
rect 3084 175 3132 333
rect 3252 234 3356 333
rect 3252 188 3281 234
rect 3327 188 3356 234
rect 3252 175 3356 188
rect 3476 175 3524 333
rect 3644 320 3732 333
rect 3644 274 3673 320
rect 3719 274 3732 320
rect 3644 175 3732 274
rect 3804 222 3892 333
rect 3804 82 3817 222
rect 3863 82 3892 222
rect 3804 69 3892 82
rect 4012 320 4116 333
rect 4012 180 4041 320
rect 4087 180 4116 320
rect 4012 69 4116 180
rect 4236 222 4340 333
rect 4236 82 4265 222
rect 4311 82 4340 222
rect 4236 69 4340 82
rect 4460 320 4564 333
rect 4460 180 4489 320
rect 4535 180 4564 320
rect 4460 69 4564 180
rect 4684 222 4772 333
rect 4684 82 4713 222
rect 4759 82 4772 222
rect 4684 69 4772 82
<< mvpdiff >>
rect 1448 955 1520 968
rect 36 739 124 849
rect 36 599 49 739
rect 95 599 124 739
rect 36 573 124 599
rect 224 836 328 849
rect 224 696 253 836
rect 299 696 328 836
rect 224 573 328 696
rect 428 726 516 849
rect 1448 909 1461 955
rect 1507 909 1520 955
rect 2088 955 2160 968
rect 1448 890 1520 909
rect 2088 909 2101 955
rect 2147 909 2160 955
rect 2088 896 2160 909
rect 2088 890 2148 896
rect 1448 773 1580 890
rect 428 586 457 726
rect 503 586 516 726
rect 428 573 516 586
rect 588 760 676 773
rect 588 714 601 760
rect 647 714 676 760
rect 588 573 676 714
rect 776 726 880 773
rect 776 586 805 726
rect 851 586 880 726
rect 776 573 880 586
rect 980 726 1084 773
rect 980 586 1009 726
rect 1055 586 1084 726
rect 980 573 1084 586
rect 1184 727 1288 773
rect 1184 681 1213 727
rect 1259 681 1288 727
rect 1184 573 1288 681
rect 1388 690 1580 773
rect 1680 749 1768 890
rect 1680 703 1709 749
rect 1755 703 1768 749
rect 1680 690 1768 703
rect 1840 749 1928 890
rect 1840 703 1853 749
rect 1899 703 1928 749
rect 1840 690 1928 703
rect 2028 773 2148 890
rect 3836 926 3924 939
rect 2876 836 2964 849
rect 2876 790 2889 836
rect 2935 790 2964 836
rect 2028 690 2208 773
rect 1388 573 1468 690
rect 2128 573 2208 690
rect 2308 726 2412 773
rect 2308 586 2337 726
rect 2383 586 2412 726
rect 2308 573 2412 586
rect 2512 726 2616 773
rect 2512 586 2541 726
rect 2587 586 2616 726
rect 2512 573 2616 586
rect 2716 632 2804 773
rect 2716 586 2745 632
rect 2791 586 2804 632
rect 2716 573 2804 586
rect 2876 573 2964 790
rect 3064 632 3168 849
rect 3064 586 3093 632
rect 3139 586 3168 632
rect 3064 573 3168 586
rect 3268 836 3372 849
rect 3268 790 3297 836
rect 3343 790 3372 836
rect 3268 573 3372 790
rect 3472 632 3576 849
rect 3472 586 3501 632
rect 3547 586 3576 632
rect 3472 573 3576 586
rect 3676 836 3764 849
rect 3676 696 3705 836
rect 3751 696 3764 836
rect 3676 573 3764 696
rect 3836 786 3849 926
rect 3895 786 3924 926
rect 3836 573 3924 786
rect 4024 726 4128 939
rect 4024 586 4053 726
rect 4099 586 4128 726
rect 4024 573 4128 586
rect 4228 926 4332 939
rect 4228 786 4257 926
rect 4303 786 4332 926
rect 4228 573 4332 786
rect 4432 726 4536 939
rect 4432 586 4461 726
rect 4507 586 4536 726
rect 4432 573 4536 586
rect 4636 926 4724 939
rect 4636 786 4665 926
rect 4711 786 4724 926
rect 4636 573 4724 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 657 228 703 274
rect 881 274 927 320
rect 1105 274 1151 320
rect 1729 228 1775 274
rect 2121 274 2167 320
rect 2345 274 2391 320
rect 2569 273 2615 319
rect 2889 251 2935 297
rect 3281 188 3327 234
rect 3673 274 3719 320
rect 3817 82 3863 222
rect 4041 180 4087 320
rect 4265 82 4311 222
rect 4489 180 4535 320
rect 4713 82 4759 222
<< mvpdiffc >>
rect 49 599 95 739
rect 253 696 299 836
rect 1461 909 1507 955
rect 2101 909 2147 955
rect 457 586 503 726
rect 601 714 647 760
rect 805 586 851 726
rect 1009 586 1055 726
rect 1213 681 1259 727
rect 1709 703 1755 749
rect 1853 703 1899 749
rect 2889 790 2935 836
rect 2337 586 2383 726
rect 2541 586 2587 726
rect 2745 586 2791 632
rect 3093 586 3139 632
rect 3297 790 3343 836
rect 3501 586 3547 632
rect 3705 696 3751 836
rect 3849 786 3895 926
rect 4053 586 4099 726
rect 4257 786 4303 926
rect 4461 586 4507 726
rect 4665 786 4711 926
<< polysilicon >>
rect 328 913 1184 953
rect 124 849 224 893
rect 328 849 428 913
rect 880 852 980 865
rect 676 773 776 817
rect 880 806 921 852
rect 967 806 980 852
rect 880 773 980 806
rect 1084 852 1184 913
rect 1084 806 1125 852
rect 1171 806 1184 852
rect 1580 890 1680 934
rect 1928 890 2028 934
rect 2268 913 3064 953
rect 3924 939 4024 983
rect 4128 939 4228 983
rect 4332 939 4432 983
rect 4536 939 4636 983
rect 1084 773 1184 806
rect 1288 773 1388 817
rect 2268 843 2308 913
rect 2208 773 2308 843
rect 2412 852 2512 865
rect 2412 806 2453 852
rect 2499 806 2512 852
rect 2964 849 3064 913
rect 3168 849 3268 893
rect 3372 849 3472 893
rect 3576 849 3676 893
rect 2412 773 2512 806
rect 2616 773 2716 817
rect 124 497 224 573
rect 328 529 428 573
rect 676 529 776 573
rect 124 451 137 497
rect 183 451 224 497
rect 124 377 224 451
rect 348 412 428 529
rect 124 333 244 377
rect 348 366 361 412
rect 407 377 428 412
rect 732 513 776 529
rect 732 500 804 513
rect 732 454 745 500
rect 791 454 804 500
rect 732 377 804 454
rect 880 465 980 573
rect 1084 529 1184 573
rect 1288 529 1388 573
rect 1348 493 1388 529
rect 1348 480 1468 493
rect 880 425 1300 465
rect 1180 412 1300 425
rect 407 366 468 377
rect 348 333 468 366
rect 732 333 852 377
rect 956 333 1076 377
rect 1180 366 1197 412
rect 1243 366 1300 412
rect 1180 333 1300 366
rect 1348 434 1361 480
rect 1407 434 1468 480
rect 1348 333 1468 434
rect 1580 377 1680 690
rect 1928 585 2028 690
rect 1852 572 2028 585
rect 1852 526 1865 572
rect 1911 545 2028 572
rect 1911 526 1924 545
rect 1852 377 1924 526
rect 2208 465 2308 573
rect 2412 529 2512 573
rect 2616 529 2716 573
rect 1580 333 1700 377
rect 1804 333 1924 377
rect 1972 425 2308 465
rect 1972 333 2092 425
rect 2420 377 2512 529
rect 2676 398 2716 529
rect 2964 412 3064 573
rect 2196 333 2316 377
rect 2420 333 2540 377
rect 2676 369 2760 398
rect 124 131 244 175
rect 348 115 468 175
rect 732 171 852 215
rect 956 115 1076 215
rect 1180 171 1300 215
rect 1348 171 1468 215
rect 348 75 1076 115
rect 1580 75 1700 215
rect 1804 171 1924 215
rect 1972 171 2092 215
rect 2196 182 2316 215
rect 2196 136 2209 182
rect 2255 136 2316 182
rect 2420 171 2540 215
rect 2688 182 2760 369
rect 2964 366 2977 412
rect 3023 377 3064 412
rect 3168 529 3268 573
rect 3372 531 3472 573
rect 3168 420 3252 529
rect 3168 377 3193 420
rect 3023 366 3084 377
rect 2964 333 3084 366
rect 3132 374 3193 377
rect 3239 374 3252 420
rect 3372 485 3409 531
rect 3455 485 3472 531
rect 3372 377 3472 485
rect 3576 540 3676 573
rect 3576 494 3593 540
rect 3639 494 3676 540
rect 3576 482 3676 494
rect 3576 377 3644 482
rect 3924 465 4024 573
rect 4128 465 4228 573
rect 4332 465 4432 573
rect 4536 465 4636 573
rect 3132 333 3252 374
rect 3356 333 3476 377
rect 3524 333 3644 377
rect 3892 452 4684 465
rect 3892 406 3905 452
rect 3951 406 4155 452
rect 4201 406 4368 452
rect 4414 406 4684 452
rect 3892 393 4684 406
rect 3892 333 4012 393
rect 4116 333 4236 393
rect 4340 333 4460 393
rect 4564 333 4684 393
rect 2196 123 2316 136
rect 2688 136 2701 182
rect 2747 136 2760 182
rect 2688 123 2760 136
rect 2964 131 3084 175
rect 3132 131 3252 175
rect 3356 75 3476 175
rect 3524 131 3644 175
rect 1580 35 3476 75
rect 3892 25 4012 69
rect 4116 25 4236 69
rect 4340 25 4460 69
rect 4564 25 4684 69
<< polycontact >>
rect 921 806 967 852
rect 1125 806 1171 852
rect 2453 806 2499 852
rect 137 451 183 497
rect 361 366 407 412
rect 745 454 791 500
rect 1197 366 1243 412
rect 1361 434 1407 480
rect 1865 526 1911 572
rect 2209 136 2255 182
rect 2977 366 3023 412
rect 3193 374 3239 420
rect 3409 485 3455 531
rect 3593 494 3639 540
rect 3905 406 3951 452
rect 4155 406 4201 452
rect 4368 406 4414 452
rect 2701 136 2747 182
<< metal1 >>
rect 0 955 4816 1098
rect 0 918 1461 955
rect 253 836 299 918
rect 49 739 95 750
rect 601 760 647 918
rect 1507 918 2101 955
rect 1461 898 1507 909
rect 2147 926 4816 955
rect 2147 918 3849 926
rect 2101 898 2147 909
rect 253 685 299 696
rect 457 726 503 737
rect 95 599 407 634
rect 49 588 407 599
rect 137 497 315 542
rect 183 451 315 497
rect 137 440 315 451
rect 361 412 407 588
rect 361 348 407 366
rect 49 320 407 348
rect 95 302 407 320
rect 601 703 647 714
rect 693 852 967 863
rect 693 806 921 852
rect 1114 806 1125 852
rect 1171 806 2453 852
rect 2499 806 2510 852
rect 2878 836 2946 918
rect 693 795 967 806
rect 693 657 739 795
rect 2878 790 2889 836
rect 2935 790 2946 836
rect 3286 836 3354 918
rect 3286 790 3297 836
rect 3343 790 3354 836
rect 3705 836 3751 918
rect 1213 749 1755 760
rect 503 611 739 657
rect 805 726 851 737
rect 503 586 543 611
rect 457 320 543 586
rect 1009 726 1055 737
rect 851 586 927 592
rect 805 546 927 586
rect 1213 727 1709 749
rect 1259 703 1709 727
rect 1259 681 1755 703
rect 1853 749 2383 760
rect 1899 726 2383 749
rect 1899 714 2337 726
rect 1899 703 2167 714
rect 1853 692 2167 703
rect 1213 670 1755 681
rect 1055 586 1911 621
rect 1009 575 1911 586
rect 589 500 754 542
rect 589 454 745 500
rect 791 454 802 500
rect 49 263 95 274
rect 457 274 497 320
rect 881 320 927 546
rect 457 263 543 274
rect 657 274 703 285
rect 273 234 319 245
rect 273 90 319 188
rect 881 263 927 274
rect 1105 320 1151 575
rect 1865 572 1911 575
rect 1865 515 1911 526
rect 1361 480 1407 491
rect 2121 469 2167 692
rect 2337 575 2383 586
rect 2541 726 3639 737
rect 2587 691 3639 726
rect 1407 434 2167 469
rect 1361 423 2167 434
rect 1197 412 1243 423
rect 1243 366 2075 377
rect 1197 331 2075 366
rect 1105 263 1151 274
rect 1729 274 1775 285
rect 657 90 703 228
rect 1729 90 1775 228
rect 2029 182 2075 331
rect 2121 320 2167 423
rect 2541 422 2587 586
rect 2121 263 2167 274
rect 2345 376 2587 422
rect 2745 632 2791 643
rect 2345 320 2391 376
rect 2745 330 2791 586
rect 3090 632 3139 643
rect 3090 586 3093 632
rect 3090 575 3139 586
rect 3501 632 3547 643
rect 2852 412 3023 430
rect 2852 366 2977 412
rect 2852 354 3023 366
rect 2345 263 2391 274
rect 2569 319 2791 330
rect 2615 308 2791 319
rect 3090 308 3136 575
rect 3237 531 3455 542
rect 3237 485 3409 531
rect 3237 466 3455 485
rect 3501 423 3547 586
rect 3593 540 3639 691
rect 3895 918 4257 926
rect 3849 775 3895 786
rect 4303 918 4665 926
rect 4257 775 4303 786
rect 4711 918 4816 926
rect 4665 775 4711 786
rect 3705 685 3751 696
rect 4041 726 4099 737
rect 4041 586 4053 726
rect 4461 726 4577 737
rect 4099 586 4461 621
rect 4507 586 4577 726
rect 4041 575 4577 586
rect 3593 483 3639 494
rect 3904 452 4414 463
rect 3904 423 3905 452
rect 3501 420 3905 423
rect 3182 374 3193 420
rect 3239 406 3905 420
rect 3951 406 4155 452
rect 4201 406 4368 452
rect 3239 395 4414 406
rect 3239 374 3951 395
rect 2615 297 3136 308
rect 2615 273 2889 297
rect 2569 251 2889 273
rect 2935 251 3136 297
rect 3673 373 3951 374
rect 3673 320 3719 373
rect 4460 331 4577 575
rect 3673 263 3719 274
rect 4041 320 4577 331
rect 2569 240 3136 251
rect 3281 234 3327 245
rect 2029 136 2209 182
rect 2255 136 2701 182
rect 2747 136 2758 182
rect 3281 90 3327 188
rect 3817 222 3863 233
rect 0 82 3817 90
rect 4087 279 4489 320
rect 4041 169 4087 180
rect 4265 222 4311 233
rect 3863 82 4265 90
rect 4535 180 4577 320
rect 4489 169 4577 180
rect 4713 222 4759 233
rect 4311 82 4713 90
rect 4759 82 4816 90
rect 0 -90 4816 82
<< labels >>
flabel metal1 s 137 440 315 542 0 FreeSans 200 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 589 500 754 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4461 621 4577 737 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3237 466 3455 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 2852 354 3023 430 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 918 4816 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 1729 245 1775 285 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 589 454 802 500 1 D
port 1 nsew default input
rlabel metal1 s 4041 621 4099 737 1 Q
port 5 nsew default output
rlabel metal1 s 4041 575 4577 621 1 Q
port 5 nsew default output
rlabel metal1 s 4460 331 4577 575 1 Q
port 5 nsew default output
rlabel metal1 s 4041 279 4577 331 1 Q
port 5 nsew default output
rlabel metal1 s 4489 169 4577 279 1 Q
port 5 nsew default output
rlabel metal1 s 4041 169 4087 279 1 Q
port 5 nsew default output
rlabel metal1 s 4665 898 4711 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4257 898 4303 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3849 898 3895 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3705 898 3751 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3286 898 3354 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2878 898 2946 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2101 898 2147 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1461 898 1507 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 898 647 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 898 299 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4665 790 4711 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4257 790 4303 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3849 790 3895 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3705 790 3751 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3286 790 3354 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2878 790 2946 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 790 647 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 790 299 898 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4665 775 4711 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4257 775 4303 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3849 775 3895 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3705 775 3751 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 775 647 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 775 299 790 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3705 703 3751 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 601 703 647 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 703 299 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3705 685 3751 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 253 685 299 703 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 657 245 703 285 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3281 233 3327 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1729 233 1775 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 657 233 703 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 233 319 245 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4713 90 4759 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4265 90 4311 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3817 90 3863 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3281 90 3327 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1729 90 1775 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 657 90 703 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4816 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 1008
string GDS_END 652202
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 641190
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
