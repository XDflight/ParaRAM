magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 3808 844
rect 69 496 115 724
rect 466 430 542 654
rect 1256 521 1302 724
rect 58 354 318 430
rect 373 354 542 430
rect 1938 584 1984 724
rect 262 60 330 199
rect 1213 60 1281 215
rect 2327 552 2373 724
rect 2740 608 2786 724
rect 2940 542 2995 639
rect 3148 608 3194 724
rect 3352 542 3398 639
rect 3556 609 3602 724
rect 2940 466 3678 542
rect 2021 318 2213 353
rect 2021 307 2551 318
rect 3602 307 3678 466
rect 2157 242 2551 307
rect 2964 253 3678 307
rect 1964 60 2010 169
rect 2740 60 2786 161
rect 2964 141 3010 253
rect 3188 60 3234 161
rect 3412 141 3458 253
rect 3636 60 3682 161
rect 0 -60 3808 60
<< obsm1 >>
rect 762 512 808 625
rect 1464 632 1879 678
rect 600 466 1087 512
rect 38 245 423 292
rect 38 153 106 245
rect 377 199 423 245
rect 600 199 646 466
rect 692 374 987 420
rect 692 289 738 374
rect 1041 315 1087 466
rect 1464 407 1510 632
rect 1729 407 1786 570
rect 1833 538 1879 632
rect 2040 632 2281 678
rect 2040 538 2086 632
rect 1833 491 2086 538
rect 2143 445 2189 570
rect 1137 361 1510 407
rect 1041 268 1416 315
rect 377 153 554 199
rect 600 153 778 199
rect 1464 156 1510 361
rect 1583 361 1786 407
rect 1835 399 2189 445
rect 2235 445 2281 632
rect 2536 537 2582 653
rect 2536 491 2786 537
rect 2235 399 2683 445
rect 1583 152 1655 361
rect 1835 261 1883 399
rect 2615 393 2683 399
rect 2740 419 2786 491
rect 2740 365 3514 419
rect 2740 307 2786 365
rect 1835 215 2102 261
rect 2621 253 2786 307
rect 1583 106 1815 152
rect 2056 152 2102 215
rect 2621 152 2667 253
rect 2056 106 2247 152
rect 2319 106 2667 152
<< labels >>
rlabel metal1 s 2021 318 2213 353 6 CLK
port 1 nsew clock input
rlabel metal1 s 2021 307 2551 318 6 CLK
port 1 nsew clock input
rlabel metal1 s 2157 242 2551 307 6 CLK
port 1 nsew clock input
rlabel metal1 s 466 430 542 654 6 E
port 2 nsew default input
rlabel metal1 s 373 354 542 430 6 E
port 2 nsew default input
rlabel metal1 s 58 354 318 430 6 TE
port 3 nsew default input
rlabel metal1 s 3352 542 3398 639 6 Q
port 4 nsew default output
rlabel metal1 s 2940 542 2995 639 6 Q
port 4 nsew default output
rlabel metal1 s 2940 466 3678 542 6 Q
port 4 nsew default output
rlabel metal1 s 3602 307 3678 466 6 Q
port 4 nsew default output
rlabel metal1 s 2964 253 3678 307 6 Q
port 4 nsew default output
rlabel metal1 s 3412 141 3458 253 6 Q
port 4 nsew default output
rlabel metal1 s 2964 141 3010 253 6 Q
port 4 nsew default output
rlabel metal1 s 0 724 3808 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3556 609 3602 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3148 609 3194 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 609 2786 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 609 2373 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 609 1984 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 609 1302 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 609 115 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3148 608 3194 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 608 2786 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 608 2373 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 608 1984 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 608 1302 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 608 115 609 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 584 2373 608 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 584 1984 608 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 584 1302 608 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 584 115 608 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 552 2373 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 552 1302 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 552 115 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1256 521 1302 552 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 521 115 552 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 521 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1213 199 1281 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 169 1281 199 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 169 330 199 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1964 161 2010 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 161 1281 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 161 330 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3636 60 3682 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3188 60 3234 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2740 60 2786 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1964 60 2010 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 465242
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 457096
<< end >>
