magic
tech gf180mcuC
timestamp 1667403419
<< metal1 >>
rect 0 111 62 123
rect 11 70 16 111
rect 28 76 33 104
rect 26 70 36 76
rect 45 70 50 111
rect 12 44 22 50
rect 28 35 33 70
rect 40 57 50 63
rect 14 30 33 35
rect 14 19 19 30
rect 42 12 47 36
rect 0 0 62 12
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 9 112 19 118
rect 33 112 43 118
rect 10 111 18 112
rect 34 111 42 112
rect 26 69 36 77
rect 40 56 50 64
rect 12 43 22 51
rect 10 11 18 12
rect 34 11 42 12
rect 9 5 19 11
rect 33 5 43 11
rect 10 4 18 5
rect 34 4 42 5
<< labels >>
rlabel metal2 s 12 43 22 51 6 A
port 1 nsew signal input
rlabel metal1 s 12 44 22 50 6 A
port 1 nsew signal input
rlabel metal2 s 40 56 50 64 6 B
port 2 nsew signal input
rlabel metal1 s 40 57 50 63 6 B
port 2 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 45 70 50 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 111 62 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 42 0 47 36 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 62 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 26 69 36 77 6 Y
port 5 nsew signal output
rlabel metal1 s 14 19 19 35 6 Y
port 5 nsew signal output
rlabel metal1 s 14 30 33 35 6 Y
port 5 nsew signal output
rlabel metal1 s 28 30 33 104 6 Y
port 5 nsew signal output
rlabel metal1 s 26 70 36 76 6 Y
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 62 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
