magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 5238 1094
<< pwell >>
rect -86 -86 5238 453
<< mvnmos >>
rect 129 157 249 275
rect 353 157 473 275
rect 521 157 641 275
rect 745 157 865 275
rect 913 157 1033 275
rect 1328 157 1448 315
rect 1552 157 1672 315
rect 1920 215 2040 333
rect 2144 215 2264 333
rect 2312 215 2432 333
rect 2536 215 2656 333
rect 2864 215 2984 333
rect 3032 215 3152 333
rect 3256 215 3376 333
rect 3480 215 3600 333
rect 3888 157 4008 275
rect 4056 157 4176 275
rect 4280 157 4400 275
rect 4540 157 4660 315
rect 4908 69 5028 333
<< mvpmos >>
rect 139 651 239 851
rect 343 651 443 851
rect 491 651 591 851
rect 745 651 845 851
rect 893 651 993 851
rect 1288 584 1388 860
rect 1492 584 1592 860
rect 1844 591 1944 791
rect 2048 591 2148 791
rect 2252 591 2352 791
rect 2536 591 2636 791
rect 2884 626 2984 826
rect 3168 592 3268 792
rect 3372 592 3472 792
rect 3576 592 3676 792
rect 3930 684 4030 884
rect 4134 684 4234 884
rect 4382 636 4482 912
rect 4586 636 4686 912
rect 4826 573 4926 939
<< mvndiff >>
rect 1240 302 1328 315
rect 41 216 129 275
rect 41 170 54 216
rect 100 170 129 216
rect 41 157 129 170
rect 249 216 353 275
rect 249 170 278 216
rect 324 170 353 216
rect 249 157 353 170
rect 473 157 521 275
rect 641 216 745 275
rect 641 170 670 216
rect 716 170 745 216
rect 641 157 745 170
rect 865 157 913 275
rect 1033 157 1165 275
rect 1240 256 1253 302
rect 1299 256 1328 302
rect 1240 157 1328 256
rect 1448 216 1552 315
rect 1448 170 1477 216
rect 1523 170 1552 216
rect 1448 157 1552 170
rect 1672 302 1760 315
rect 1672 256 1701 302
rect 1747 256 1760 302
rect 1672 157 1760 256
rect 1832 274 1920 333
rect 1832 228 1845 274
rect 1891 228 1920 274
rect 1832 215 1920 228
rect 2040 274 2144 333
rect 2040 228 2069 274
rect 2115 228 2144 274
rect 2040 215 2144 228
rect 2264 215 2312 333
rect 2432 215 2536 333
rect 2656 274 2864 333
rect 2656 228 2685 274
rect 2731 228 2864 274
rect 2656 215 2864 228
rect 2984 215 3032 333
rect 3152 320 3256 333
rect 3152 274 3181 320
rect 3227 274 3256 320
rect 3152 215 3256 274
rect 3376 320 3480 333
rect 3376 274 3405 320
rect 3451 274 3480 320
rect 3376 215 3480 274
rect 3600 320 3688 333
rect 3600 274 3629 320
rect 3675 274 3688 320
rect 4460 275 4540 315
rect 3600 215 3688 274
rect 3800 216 3888 275
rect 1093 96 1165 157
rect 1093 50 1106 96
rect 1152 50 1165 96
rect 1093 37 1165 50
rect 3800 170 3813 216
rect 3859 170 3888 216
rect 3800 157 3888 170
rect 4008 157 4056 275
rect 4176 216 4280 275
rect 4176 170 4205 216
rect 4251 170 4280 216
rect 4176 157 4280 170
rect 4400 157 4540 275
rect 4660 216 4748 315
rect 4660 170 4689 216
rect 4735 170 4748 216
rect 4660 157 4748 170
rect 4820 309 4908 333
rect 4820 169 4833 309
rect 4879 169 4908 309
rect 4820 69 4908 169
rect 5028 320 5116 333
rect 5028 180 5057 320
rect 5103 180 5116 320
rect 5028 69 5116 180
<< mvpdiff >>
rect 3036 958 3108 971
rect 51 804 139 851
rect 51 664 64 804
rect 110 664 139 804
rect 51 651 139 664
rect 239 838 343 851
rect 239 698 268 838
rect 314 698 343 838
rect 239 651 343 698
rect 443 651 491 851
rect 591 838 745 851
rect 591 698 670 838
rect 716 698 745 838
rect 591 651 745 698
rect 845 651 893 851
rect 993 838 1081 851
rect 993 792 1022 838
rect 1068 792 1081 838
rect 993 651 1081 792
rect 1200 645 1288 860
rect 1200 599 1213 645
rect 1259 599 1288 645
rect 1200 584 1288 599
rect 1388 847 1492 860
rect 1388 801 1417 847
rect 1463 801 1492 847
rect 1388 584 1492 801
rect 1592 643 1680 860
rect 2412 923 2484 936
rect 2412 877 2425 923
rect 2471 877 2484 923
rect 3036 912 3049 958
rect 3095 912 3108 958
rect 3036 900 3108 912
rect 2412 865 2484 877
rect 2412 791 2476 865
rect 3044 826 3108 900
rect 1592 597 1621 643
rect 1667 597 1680 643
rect 1592 584 1680 597
rect 1756 744 1844 791
rect 1756 604 1769 744
rect 1815 604 1844 744
rect 1756 591 1844 604
rect 1944 778 2048 791
rect 1944 638 1973 778
rect 2019 638 2048 778
rect 1944 591 2048 638
rect 2148 710 2252 791
rect 2148 664 2177 710
rect 2223 664 2252 710
rect 2148 591 2252 664
rect 2352 591 2536 791
rect 2636 710 2724 791
rect 2636 664 2665 710
rect 2711 664 2724 710
rect 2636 591 2724 664
rect 2796 710 2884 826
rect 2796 664 2809 710
rect 2855 664 2884 710
rect 2796 626 2884 664
rect 2984 792 3108 826
rect 4746 912 4826 939
rect 4294 899 4382 912
rect 4294 884 4307 899
rect 3842 871 3930 884
rect 3842 825 3855 871
rect 3901 825 3930 871
rect 2984 626 3168 792
rect 3088 592 3168 626
rect 3268 768 3372 792
rect 3268 628 3297 768
rect 3343 628 3372 768
rect 3268 592 3372 628
rect 3472 779 3576 792
rect 3472 639 3501 779
rect 3547 639 3576 779
rect 3472 592 3576 639
rect 3676 651 3764 792
rect 3842 684 3930 825
rect 4030 743 4134 884
rect 4030 697 4059 743
rect 4105 697 4134 743
rect 4030 684 4134 697
rect 4234 853 4307 884
rect 4353 853 4382 899
rect 4234 684 4382 853
rect 3676 605 3705 651
rect 3751 605 3764 651
rect 3676 592 3764 605
rect 4302 636 4382 684
rect 4482 695 4586 912
rect 4482 649 4511 695
rect 4557 649 4586 695
rect 4482 636 4586 649
rect 4686 899 4826 912
rect 4686 759 4715 899
rect 4761 759 4826 899
rect 4686 636 4826 759
rect 4746 573 4826 636
rect 4926 804 5014 939
rect 4926 664 4955 804
rect 5001 664 5014 804
rect 4926 573 5014 664
<< mvndiffc >>
rect 54 170 100 216
rect 278 170 324 216
rect 670 170 716 216
rect 1253 256 1299 302
rect 1477 170 1523 216
rect 1701 256 1747 302
rect 1845 228 1891 274
rect 2069 228 2115 274
rect 2685 228 2731 274
rect 3181 274 3227 320
rect 3405 274 3451 320
rect 3629 274 3675 320
rect 1106 50 1152 96
rect 3813 170 3859 216
rect 4205 170 4251 216
rect 4689 170 4735 216
rect 4833 169 4879 309
rect 5057 180 5103 320
<< mvpdiffc >>
rect 64 664 110 804
rect 268 698 314 838
rect 670 698 716 838
rect 1022 792 1068 838
rect 1213 599 1259 645
rect 1417 801 1463 847
rect 2425 877 2471 923
rect 3049 912 3095 958
rect 1621 597 1667 643
rect 1769 604 1815 744
rect 1973 638 2019 778
rect 2177 664 2223 710
rect 2665 664 2711 710
rect 2809 664 2855 710
rect 3855 825 3901 871
rect 3297 628 3343 768
rect 3501 639 3547 779
rect 4059 697 4105 743
rect 4307 853 4353 899
rect 3705 605 3751 651
rect 4511 649 4557 695
rect 4715 759 4761 899
rect 4955 664 5001 804
<< polysilicon >>
rect 139 943 993 983
rect 139 851 239 943
rect 343 851 443 895
rect 491 851 591 895
rect 745 851 845 895
rect 893 851 993 943
rect 1492 943 2148 983
rect 1288 860 1388 904
rect 1492 860 1592 943
rect 2048 870 2148 943
rect 139 499 239 651
rect 343 607 443 651
rect 129 486 239 499
rect 129 440 142 486
rect 188 440 239 486
rect 129 319 239 440
rect 353 486 425 607
rect 491 499 591 651
rect 353 440 366 486
rect 412 440 425 486
rect 353 319 425 440
rect 485 486 591 499
rect 485 440 498 486
rect 544 440 591 486
rect 485 427 591 440
rect 745 486 845 651
rect 893 607 993 651
rect 1844 791 1944 835
rect 2048 824 2089 870
rect 2135 824 2148 870
rect 2048 791 2148 824
rect 2252 791 2352 835
rect 2536 791 2636 835
rect 2884 826 2984 870
rect 3168 944 4030 984
rect 3168 792 3268 944
rect 3930 884 4030 944
rect 4134 884 4234 928
rect 4382 912 4482 956
rect 4586 912 4686 956
rect 4826 939 4926 983
rect 3372 871 3472 884
rect 3372 825 3385 871
rect 3431 825 3472 871
rect 3372 792 3472 825
rect 3576 792 3676 836
rect 1288 542 1388 584
rect 745 440 758 486
rect 804 440 845 486
rect 745 319 845 440
rect 913 486 1033 499
rect 913 440 946 486
rect 992 440 1033 486
rect 1288 496 1301 542
rect 1347 496 1388 542
rect 1288 483 1388 496
rect 129 275 249 319
rect 353 275 473 319
rect 521 275 641 319
rect 745 275 865 319
rect 913 275 1033 440
rect 1328 359 1388 483
rect 1492 486 1592 584
rect 1492 440 1505 486
rect 1551 440 1592 486
rect 1492 427 1592 440
rect 1844 499 1944 591
rect 2048 547 2148 591
rect 2252 547 2352 591
rect 2312 499 2352 547
rect 1844 486 2264 499
rect 1844 440 1857 486
rect 1903 440 2185 486
rect 2231 440 2264 486
rect 1844 427 2264 440
rect 1552 359 1592 427
rect 1328 315 1448 359
rect 1552 315 1672 359
rect 1920 333 2040 377
rect 2144 333 2264 427
rect 2312 486 2432 499
rect 2312 440 2373 486
rect 2419 440 2432 486
rect 2312 333 2432 440
rect 2536 377 2636 591
rect 2884 578 2984 626
rect 3930 640 4030 684
rect 2884 532 2897 578
rect 2943 532 2984 578
rect 2884 377 2984 532
rect 3168 548 3268 592
rect 3372 548 3472 592
rect 3576 548 3676 592
rect 3168 465 3208 548
rect 2536 333 2656 377
rect 2864 333 2984 377
rect 3032 393 3208 465
rect 3432 465 3472 548
rect 3636 499 3676 548
rect 3636 486 3780 499
rect 3432 393 3580 465
rect 3636 440 3721 486
rect 3767 440 3780 486
rect 3636 427 3780 440
rect 3930 486 4008 640
rect 3930 440 3949 486
rect 3995 440 4008 486
rect 3032 333 3152 393
rect 3480 377 3580 393
rect 3256 333 3376 377
rect 3480 333 3600 377
rect 3930 319 4008 440
rect 4134 486 4234 684
rect 4382 499 4482 636
rect 4134 440 4175 486
rect 4221 440 4234 486
rect 4134 394 4234 440
rect 3888 275 4008 319
rect 4056 335 4234 394
rect 4300 486 4482 499
rect 4300 440 4313 486
rect 4359 440 4482 486
rect 4300 429 4482 440
rect 4586 486 4686 636
rect 4586 440 4603 486
rect 4649 440 4686 486
rect 4586 433 4686 440
rect 4826 486 4926 573
rect 4826 440 4839 486
rect 4885 463 4926 486
rect 4885 440 5028 463
rect 4056 275 4176 335
rect 4300 319 4400 429
rect 4586 359 4660 433
rect 4826 393 5028 440
rect 4280 275 4400 319
rect 4540 315 4660 359
rect 4908 333 5028 393
rect 129 65 249 157
rect 353 113 473 157
rect 521 65 641 157
rect 745 113 865 157
rect 913 113 1033 157
rect 129 25 641 65
rect 1328 113 1448 157
rect 1552 97 1672 157
rect 1920 97 2040 215
rect 2144 171 2264 215
rect 2312 171 2432 215
rect 1552 25 2040 97
rect 2536 65 2656 215
rect 2864 171 2984 215
rect 3032 171 3152 215
rect 3256 182 3376 215
rect 3256 136 3269 182
rect 3315 136 3376 182
rect 3480 171 3600 215
rect 3256 123 3376 136
rect 3888 113 4008 157
rect 4056 113 4176 157
rect 4280 65 4400 157
rect 4540 113 4660 157
rect 2536 25 4400 65
rect 4908 25 5028 69
<< polycontact >>
rect 142 440 188 486
rect 366 440 412 486
rect 498 440 544 486
rect 2089 824 2135 870
rect 3385 825 3431 871
rect 758 440 804 486
rect 946 440 992 486
rect 1301 496 1347 542
rect 1505 440 1551 486
rect 1857 440 1903 486
rect 2185 440 2231 486
rect 2373 440 2419 486
rect 2897 532 2943 578
rect 3721 440 3767 486
rect 3949 440 3995 486
rect 4175 440 4221 486
rect 4313 440 4359 486
rect 4603 440 4649 486
rect 4839 440 4885 486
rect 3269 136 3315 182
<< metal1 >>
rect 0 958 5152 1098
rect 0 923 3049 958
rect 0 918 2425 923
rect 268 838 314 918
rect 64 804 110 815
rect 268 687 314 698
rect 670 838 716 849
rect 1022 838 1068 918
rect 1406 847 1474 918
rect 2471 918 3049 923
rect 3095 918 5152 958
rect 3049 901 3095 912
rect 1406 801 1417 847
rect 1463 801 1474 847
rect 2078 824 2089 870
rect 2135 824 2146 870
rect 2425 866 2471 877
rect 3855 871 3901 918
rect 3130 855 3385 871
rect 2078 820 2146 824
rect 3084 825 3385 855
rect 3431 825 3442 871
rect 4296 899 4364 918
rect 4296 853 4307 899
rect 4353 853 4364 899
rect 4715 899 4761 918
rect 3084 820 3165 825
rect 1022 781 1068 792
rect 1973 778 2019 789
rect 1106 744 1815 755
rect 1106 733 1769 744
rect 716 709 1769 733
rect 716 698 1146 709
rect 670 687 1146 698
rect 64 634 110 664
rect 1213 645 1551 656
rect 64 588 992 634
rect 1259 599 1551 645
rect 1213 588 1551 599
rect 30 486 188 542
rect 30 440 142 486
rect 30 429 188 440
rect 366 486 418 542
rect 412 440 418 486
rect 30 354 82 429
rect 366 354 418 440
rect 498 486 544 588
rect 498 308 544 440
rect 590 486 642 542
rect 946 486 992 588
rect 590 440 758 486
rect 804 440 815 486
rect 1262 496 1301 542
rect 1347 496 1426 542
rect 1262 466 1426 496
rect 1505 486 1551 588
rect 590 354 642 440
rect 946 429 992 440
rect 1621 643 1667 654
rect 1621 497 1667 597
rect 1769 593 1815 604
rect 2078 774 3165 820
rect 3855 814 3901 825
rect 3947 843 4139 846
rect 3947 800 4251 843
rect 3501 779 3547 790
rect 3297 768 3343 779
rect 2177 710 2711 721
rect 2223 664 2665 710
rect 2177 653 2711 664
rect 2809 710 3035 721
rect 2855 664 3035 710
rect 2809 653 3035 664
rect 1973 625 2019 638
rect 1973 589 2114 625
rect 1973 579 2943 589
rect 2069 578 2943 579
rect 2069 543 2897 578
rect 1621 486 1903 497
rect 1621 451 1857 486
rect 1505 411 1551 440
rect 1253 365 1551 411
rect 1701 440 1857 451
rect 1701 429 1903 440
rect 54 262 544 308
rect 1253 302 1299 365
rect 54 216 100 262
rect 1253 245 1299 256
rect 1345 273 1655 319
rect 670 216 716 227
rect 54 159 100 170
rect 267 170 278 216
rect 324 170 335 216
rect 267 90 335 170
rect 1345 199 1391 273
rect 716 170 1391 199
rect 670 153 1391 170
rect 1477 216 1523 227
rect 1106 96 1152 107
rect 0 50 1106 90
rect 1477 90 1523 170
rect 1609 199 1655 273
rect 1701 302 1747 429
rect 1701 245 1747 256
rect 1845 274 1891 285
rect 1845 199 1891 228
rect 2069 274 2115 543
rect 2897 521 2943 532
rect 2185 486 2231 497
rect 2185 377 2231 440
rect 2373 486 2419 497
rect 2989 475 3035 653
rect 2419 440 3227 475
rect 2373 429 3227 440
rect 2185 331 3135 377
rect 2069 217 2115 228
rect 2685 274 2731 285
rect 1609 153 1891 199
rect 2685 90 2731 228
rect 3089 182 3135 331
rect 3181 320 3227 429
rect 3297 309 3343 628
rect 3947 768 3993 800
rect 4122 798 4251 800
rect 4122 797 4649 798
rect 3547 722 3993 768
rect 4059 743 4105 754
rect 4205 752 4649 797
rect 3501 331 3547 639
rect 3705 651 3751 662
rect 3705 589 3751 605
rect 3227 274 3343 309
rect 3181 263 3343 274
rect 3405 320 3547 331
rect 3451 274 3547 320
rect 3405 263 3547 274
rect 3629 543 3859 589
rect 3629 320 3675 543
rect 3629 263 3675 274
rect 3721 486 3767 497
rect 3721 182 3767 440
rect 3089 136 3269 182
rect 3315 136 3767 182
rect 3813 308 3859 543
rect 3949 486 4002 542
rect 3995 440 4002 486
rect 3949 354 4002 440
rect 4059 308 4105 697
rect 4511 695 4557 706
rect 4286 486 4359 542
rect 3813 262 4105 308
rect 4164 440 4175 486
rect 4221 440 4232 486
rect 4164 308 4232 440
rect 4286 440 4313 486
rect 4286 354 4359 440
rect 4511 308 4557 649
rect 4603 486 4649 752
rect 4715 748 4761 759
rect 4955 804 5010 815
rect 5001 664 5010 804
rect 4955 512 5010 664
rect 4603 429 4649 440
rect 4839 486 4885 497
rect 4955 466 5103 512
rect 4839 412 4885 440
rect 4692 366 4885 412
rect 4692 308 4738 366
rect 5057 320 5103 466
rect 4164 262 4738 308
rect 3813 216 3859 262
rect 4689 216 4738 262
rect 3813 159 3859 170
rect 4194 170 4205 216
rect 4251 170 4262 216
rect 4194 90 4262 170
rect 4735 170 4738 216
rect 4689 159 4738 170
rect 4833 309 4879 320
rect 5057 169 5103 180
rect 4833 90 4879 169
rect 1152 50 5152 90
rect 0 -90 5152 50
<< labels >>
flabel metal1 s 1262 466 1426 542 0 FreeSans 200 0 0 0 CLK
port 6 nsew clock input
flabel metal1 s 590 486 642 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4955 512 5010 815 0 FreeSans 200 0 0 0 Q
port 7 nsew default output
flabel metal1 s 4286 354 4359 542 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 30 429 188 542 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 3949 354 4002 542 0 FreeSans 200 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 366 354 418 542 0 FreeSans 200 0 0 0 SI
port 5 nsew default input
flabel metal1 s 0 918 5152 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 4833 285 4879 320 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 590 440 815 486 1 D
port 1 nsew default input
rlabel metal1 s 590 354 642 440 1 D
port 1 nsew default input
rlabel metal1 s 30 354 82 429 1 SE
port 3 nsew default input
rlabel metal1 s 4955 466 5103 512 1 Q
port 7 nsew default output
rlabel metal1 s 5057 169 5103 466 1 Q
port 7 nsew default output
rlabel metal1 s 4715 901 4761 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4296 901 4364 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3855 901 3901 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3049 901 3095 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2425 901 2471 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1406 901 1474 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 901 1068 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 901 314 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 866 4761 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4296 866 4364 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3855 866 3901 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2425 866 2471 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1406 866 1474 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 866 1068 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 866 314 901 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 853 4761 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4296 853 4364 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3855 853 3901 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1406 853 1474 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 853 1068 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 853 314 866 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 814 4761 853 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3855 814 3901 853 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1406 814 1474 853 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 814 1068 853 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 814 314 853 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 801 4761 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1406 801 1474 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 801 1068 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 801 314 814 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 781 4761 801 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1022 781 1068 801 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 781 314 801 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4715 748 4761 781 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 748 314 781 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 268 687 314 748 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4833 227 4879 285 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2685 227 2731 285 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 216 4879 227 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2685 216 2731 227 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1477 216 1523 227 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 107 4879 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4194 107 4262 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2685 107 2731 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1477 107 1523 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 267 107 335 216 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4833 90 4879 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4194 90 4262 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2685 90 2731 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1477 90 1523 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1106 90 1152 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 267 90 335 107 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5152 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5152 1008
string GDS_END 371648
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 359920
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
