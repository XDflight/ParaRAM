magic
tech gf180mcuC
timestamp 1666464484
<< metal1 >>
rect 0 111 16 123
rect 0 0 16 12
<< labels >>
rlabel metal1 s 0 111 16 123 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 0 16 12 6 VSS
port 2 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 16 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
