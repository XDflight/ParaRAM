magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -1857 135 1857 176
rect -1857 83 -1818 135
rect -1766 83 -1607 135
rect -1555 83 -1397 135
rect -1345 83 -1186 135
rect -1134 83 -975 135
rect -923 83 -764 135
rect -712 83 -553 135
rect -501 83 -343 135
rect -291 83 -132 135
rect -80 83 80 135
rect 132 83 291 135
rect 343 83 501 135
rect 553 83 712 135
rect 764 83 923 135
rect 975 83 1134 135
rect 1186 83 1345 135
rect 1397 83 1555 135
rect 1607 83 1766 135
rect 1818 83 1857 135
rect -1857 -83 1857 83
rect -1857 -135 -1818 -83
rect -1766 -135 -1607 -83
rect -1555 -135 -1397 -83
rect -1345 -135 -1186 -83
rect -1134 -135 -975 -83
rect -923 -135 -764 -83
rect -712 -135 -553 -83
rect -501 -135 -343 -83
rect -291 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 291 -83
rect 343 -135 501 -83
rect 553 -135 712 -83
rect 764 -135 923 -83
rect 975 -135 1134 -83
rect 1186 -135 1345 -83
rect 1397 -135 1555 -83
rect 1607 -135 1766 -83
rect 1818 -135 1857 -83
rect -1857 -176 1857 -135
<< via1 >>
rect -1818 83 -1766 135
rect -1607 83 -1555 135
rect -1397 83 -1345 135
rect -1186 83 -1134 135
rect -975 83 -923 135
rect -764 83 -712 135
rect -553 83 -501 135
rect -343 83 -291 135
rect -132 83 -80 135
rect 80 83 132 135
rect 291 83 343 135
rect 501 83 553 135
rect 712 83 764 135
rect 923 83 975 135
rect 1134 83 1186 135
rect 1345 83 1397 135
rect 1555 83 1607 135
rect 1766 83 1818 135
rect -1818 -135 -1766 -83
rect -1607 -135 -1555 -83
rect -1397 -135 -1345 -83
rect -1186 -135 -1134 -83
rect -975 -135 -923 -83
rect -764 -135 -712 -83
rect -553 -135 -501 -83
rect -343 -135 -291 -83
rect -132 -135 -80 -83
rect 80 -135 132 -83
rect 291 -135 343 -83
rect 501 -135 553 -83
rect 712 -135 764 -83
rect 923 -135 975 -83
rect 1134 -135 1186 -83
rect 1345 -135 1397 -83
rect 1555 -135 1607 -83
rect 1766 -135 1818 -83
<< metal2 >>
rect -1857 135 1857 176
rect -1857 83 -1818 135
rect -1766 83 -1607 135
rect -1555 83 -1397 135
rect -1345 83 -1186 135
rect -1134 83 -975 135
rect -923 83 -764 135
rect -712 83 -553 135
rect -501 83 -343 135
rect -291 83 -132 135
rect -80 83 80 135
rect 132 83 291 135
rect 343 83 501 135
rect 553 83 712 135
rect 764 83 923 135
rect 975 83 1134 135
rect 1186 83 1345 135
rect 1397 83 1555 135
rect 1607 83 1766 135
rect 1818 83 1857 135
rect -1857 -83 1857 83
rect -1857 -135 -1818 -83
rect -1766 -135 -1607 -83
rect -1555 -135 -1397 -83
rect -1345 -135 -1186 -83
rect -1134 -135 -975 -83
rect -923 -135 -764 -83
rect -712 -135 -553 -83
rect -501 -135 -343 -83
rect -291 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 291 -83
rect 343 -135 501 -83
rect 553 -135 712 -83
rect 764 -135 923 -83
rect 975 -135 1134 -83
rect 1186 -135 1345 -83
rect 1397 -135 1555 -83
rect 1607 -135 1766 -83
rect 1818 -135 1857 -83
rect -1857 -175 1857 -135
<< properties >>
string GDS_END 862422
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 859986
<< end >>
