magic
tech gf180mcuC
magscale 1 5
timestamp 1667403444
<< checkpaint >>
rect 12400 12400 36500 36500
<< metal4 >>
rect 13400 25705 14900 35500
tri 14900 25705 15522 26327 sw
tri 13400 24010 15095 25705 ne
rect 15095 24010 15522 25705
tri 15522 24010 17217 25705 sw
tri 15095 21888 17217 24010 ne
tri 17217 21888 19339 24010 sw
tri 17217 19766 19339 21888 ne
tri 19339 19766 21461 21888 sw
tri 19339 17644 21461 19766 ne
tri 21461 17644 23583 19766 sw
tri 21461 15522 23583 17644 ne
tri 23583 15522 25705 17644 sw
tri 23583 13400 25705 15522 ne
tri 25705 14900 26327 15522 sw
rect 25705 13400 35500 14900
<< end >>
