magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 2360 958
<< polysilicon >>
rect -31 817 89 890
rect 193 817 313 890
rect 417 817 537 890
rect 641 817 761 890
rect 865 817 985 890
rect 1089 817 1209 890
rect 1313 817 1433 890
rect 1537 817 1657 890
rect 1761 817 1881 890
rect 1985 817 2105 890
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 641 -74 761 -1
rect 865 -74 985 -1
rect 1089 -74 1209 -1
rect 1313 -74 1433 -1
rect 1537 -74 1657 -1
rect 1761 -74 1881 -1
rect 1985 -74 2105 -1
use pmos_5p04310589983222_64x8m81  pmos_5p04310589983222_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 2344 938
<< properties >>
string GDS_END 409696
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 408230
<< end >>
