magic
tech gf180mcuC
timestamp 1666464484
<< properties >>
string GDS_END 9409490
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 9160590
<< end >>
