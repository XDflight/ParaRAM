magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 22162 -6340 22775 -1078
rect 22448 -12800 22838 -10246
rect 22671 -14848 23429 -14394
rect 22650 -15879 23535 -14848
rect 22681 -15880 23535 -15879
rect 22685 -22093 23539 -19542
rect 22554 -23170 23539 -22714
<< pwell >>
rect -68 59456 23468 59488
rect -68 -88 23468 -56
<< psubdiff >>
rect 22869 -16594 23345 -16534
rect 22869 -16640 22926 -16594
rect 22972 -16640 23084 -16594
rect 23130 -16640 23242 -16594
rect 23288 -16640 23345 -16594
rect 22869 -16700 23345 -16640
<< nsubdiff >>
rect 22814 -14599 23286 -14542
rect 22814 -14645 22869 -14599
rect 22915 -14645 23027 -14599
rect 23073 -14645 23185 -14599
rect 23231 -14645 23286 -14599
rect 22814 -14702 23286 -14645
rect 22697 -22919 22852 -22862
rect 22697 -22965 22751 -22919
rect 22797 -22965 22852 -22919
rect 22697 -23022 22852 -22965
rect 23241 -22919 23396 -22862
rect 23241 -22965 23295 -22919
rect 23341 -22965 23396 -22919
rect 23241 -23022 23396 -22965
<< psubdiffcont >>
rect 22926 -16640 22972 -16594
rect 23084 -16640 23130 -16594
rect 23242 -16640 23288 -16594
<< nsubdiffcont >>
rect 22869 -14645 22915 -14599
rect 23027 -14645 23073 -14599
rect 23185 -14645 23231 -14599
rect 22751 -22965 22797 -22919
rect 23295 -22965 23341 -22919
<< polysilicon >>
rect -257 59329 57 59348
rect -257 59189 -238 59329
rect -192 59194 57 59329
rect 23341 59265 23711 59348
rect 23341 59219 23592 59265
rect 23638 59219 23711 59265
rect 23341 59194 23711 59219
rect -192 59189 -173 59194
rect -257 59170 -173 59189
rect 23519 59101 23711 59194
rect 23519 59055 23592 59101
rect 23638 59055 23711 59101
rect 23519 59009 23711 59055
rect -257 57670 57 57806
rect -257 57530 -238 57670
rect -192 57652 57 57670
rect 23341 57705 23711 57806
rect 23341 57659 23592 57705
rect 23638 57659 23711 57705
rect 23341 57652 23711 57659
rect -192 57548 -173 57652
rect 23519 57548 23711 57652
rect -192 57530 57 57548
rect -257 57394 57 57530
rect 23341 57541 23711 57548
rect 23341 57495 23592 57541
rect 23638 57495 23711 57541
rect 23341 57394 23711 57495
rect -257 55870 57 56006
rect -257 55730 -238 55870
rect -192 55852 57 55870
rect 23341 55905 23711 56006
rect 23341 55859 23592 55905
rect 23638 55859 23711 55905
rect 23341 55852 23711 55859
rect -192 55748 -173 55852
rect 23519 55748 23711 55852
rect -192 55730 57 55748
rect -257 55594 57 55730
rect 23341 55741 23711 55748
rect 23341 55695 23592 55741
rect 23638 55695 23711 55741
rect 23341 55594 23711 55695
rect -257 54070 57 54206
rect -257 53930 -238 54070
rect -192 54052 57 54070
rect 23341 54105 23711 54206
rect 23341 54059 23592 54105
rect 23638 54059 23711 54105
rect 23341 54052 23711 54059
rect -192 53948 -173 54052
rect 23519 53948 23711 54052
rect -192 53930 57 53948
rect -257 53794 57 53930
rect 23341 53941 23711 53948
rect 23341 53895 23592 53941
rect 23638 53895 23711 53941
rect 23341 53794 23711 53895
rect -257 52270 57 52406
rect -257 52130 -238 52270
rect -192 52252 57 52270
rect 23341 52305 23711 52406
rect 23341 52259 23592 52305
rect 23638 52259 23711 52305
rect 23341 52252 23711 52259
rect -192 52148 -173 52252
rect 23519 52148 23711 52252
rect -192 52130 57 52148
rect -257 51994 57 52130
rect 23341 52141 23711 52148
rect 23341 52095 23592 52141
rect 23638 52095 23711 52141
rect 23341 51994 23711 52095
rect -257 50470 57 50606
rect -257 50330 -238 50470
rect -192 50452 57 50470
rect 23341 50505 23711 50606
rect 23341 50459 23592 50505
rect 23638 50459 23711 50505
rect 23341 50452 23711 50459
rect -192 50348 -173 50452
rect 23519 50348 23711 50452
rect -192 50330 57 50348
rect -257 50194 57 50330
rect 23341 50341 23711 50348
rect 23341 50295 23592 50341
rect 23638 50295 23711 50341
rect 23341 50194 23711 50295
rect -257 48670 57 48806
rect -257 48530 -238 48670
rect -192 48652 57 48670
rect 23341 48705 23711 48806
rect 23341 48659 23592 48705
rect 23638 48659 23711 48705
rect 23341 48652 23711 48659
rect -192 48548 -173 48652
rect 23519 48548 23711 48652
rect -192 48530 57 48548
rect -257 48394 57 48530
rect 23341 48541 23711 48548
rect 23341 48495 23592 48541
rect 23638 48495 23711 48541
rect 23341 48394 23711 48495
rect -257 46870 57 47006
rect -257 46730 -238 46870
rect -192 46852 57 46870
rect 23341 46905 23711 47006
rect 23341 46859 23592 46905
rect 23638 46859 23711 46905
rect 23341 46852 23711 46859
rect -192 46748 -173 46852
rect 23519 46748 23711 46852
rect -192 46730 57 46748
rect -257 46594 57 46730
rect 23341 46741 23711 46748
rect 23341 46695 23592 46741
rect 23638 46695 23711 46741
rect 23341 46594 23711 46695
rect -257 45070 57 45206
rect -257 44930 -238 45070
rect -192 45052 57 45070
rect 23341 45105 23711 45206
rect 23341 45059 23592 45105
rect 23638 45059 23711 45105
rect 23341 45052 23711 45059
rect -192 44948 -173 45052
rect 23519 44948 23711 45052
rect -192 44930 57 44948
rect -257 44794 57 44930
rect 23341 44941 23711 44948
rect 23341 44895 23592 44941
rect 23638 44895 23711 44941
rect 23341 44794 23711 44895
rect -257 43270 57 43406
rect -257 43130 -238 43270
rect -192 43252 57 43270
rect 23341 43305 23711 43406
rect 23341 43259 23592 43305
rect 23638 43259 23711 43305
rect 23341 43252 23711 43259
rect -192 43148 -173 43252
rect 23519 43148 23711 43252
rect -192 43130 57 43148
rect -257 42994 57 43130
rect 23341 43141 23711 43148
rect 23341 43095 23592 43141
rect 23638 43095 23711 43141
rect 23341 42994 23711 43095
rect -257 41470 57 41606
rect -257 41330 -238 41470
rect -192 41452 57 41470
rect 23341 41505 23711 41606
rect 23341 41459 23592 41505
rect 23638 41459 23711 41505
rect 23341 41452 23711 41459
rect -192 41348 -173 41452
rect 23519 41348 23711 41452
rect -192 41330 57 41348
rect -257 41194 57 41330
rect 23341 41341 23711 41348
rect 23341 41295 23592 41341
rect 23638 41295 23711 41341
rect 23341 41194 23711 41295
rect -257 39670 57 39806
rect -257 39530 -238 39670
rect -192 39652 57 39670
rect 23341 39705 23711 39806
rect 23341 39659 23592 39705
rect 23638 39659 23711 39705
rect 23341 39652 23711 39659
rect -192 39548 -173 39652
rect 23519 39548 23711 39652
rect -192 39530 57 39548
rect -257 39394 57 39530
rect 23341 39541 23711 39548
rect 23341 39495 23592 39541
rect 23638 39495 23711 39541
rect 23341 39394 23711 39495
rect -257 37870 57 38006
rect -257 37730 -238 37870
rect -192 37852 57 37870
rect 23341 37905 23711 38006
rect 23341 37859 23592 37905
rect 23638 37859 23711 37905
rect 23341 37852 23711 37859
rect -192 37748 -173 37852
rect 23519 37748 23711 37852
rect -192 37730 57 37748
rect -257 37594 57 37730
rect 23341 37741 23711 37748
rect 23341 37695 23592 37741
rect 23638 37695 23711 37741
rect 23341 37594 23711 37695
rect -257 36070 57 36206
rect -257 35930 -238 36070
rect -192 36052 57 36070
rect 23341 36105 23711 36206
rect 23341 36059 23592 36105
rect 23638 36059 23711 36105
rect 23341 36052 23711 36059
rect -192 35948 -173 36052
rect 23519 35948 23711 36052
rect -192 35930 57 35948
rect -257 35794 57 35930
rect 23341 35941 23711 35948
rect 23341 35895 23592 35941
rect 23638 35895 23711 35941
rect 23341 35794 23711 35895
rect -257 34270 57 34406
rect -257 34130 -238 34270
rect -192 34252 57 34270
rect 23341 34305 23711 34406
rect 23341 34259 23592 34305
rect 23638 34259 23711 34305
rect 23341 34252 23711 34259
rect -192 34148 -173 34252
rect 23519 34148 23711 34252
rect -192 34130 57 34148
rect -257 33994 57 34130
rect 23341 34141 23711 34148
rect 23341 34095 23592 34141
rect 23638 34095 23711 34141
rect 23341 33994 23711 34095
rect -257 32470 57 32606
rect -257 32330 -238 32470
rect -192 32452 57 32470
rect 23341 32505 23711 32606
rect 23341 32459 23592 32505
rect 23638 32459 23711 32505
rect 23341 32452 23711 32459
rect -192 32348 -173 32452
rect 23519 32348 23711 32452
rect -192 32330 57 32348
rect -257 32194 57 32330
rect 23341 32341 23711 32348
rect 23341 32295 23592 32341
rect 23638 32295 23711 32341
rect 23341 32194 23711 32295
rect -257 30670 57 30806
rect -257 30530 -238 30670
rect -192 30652 57 30670
rect 23341 30705 23711 30806
rect 23341 30659 23592 30705
rect 23638 30659 23711 30705
rect 23341 30652 23711 30659
rect -192 30548 -173 30652
rect 23519 30548 23711 30652
rect -192 30530 57 30548
rect -257 30394 57 30530
rect 23341 30541 23711 30548
rect 23341 30495 23592 30541
rect 23638 30495 23711 30541
rect 23341 30394 23711 30495
rect -257 28870 57 29006
rect -257 28730 -238 28870
rect -192 28852 57 28870
rect 23341 28905 23711 29006
rect 23341 28859 23592 28905
rect 23638 28859 23711 28905
rect 23341 28852 23711 28859
rect -192 28748 -173 28852
rect 23519 28748 23711 28852
rect -192 28730 57 28748
rect -257 28594 57 28730
rect 23341 28741 23711 28748
rect 23341 28695 23592 28741
rect 23638 28695 23711 28741
rect 23341 28594 23711 28695
rect -257 27070 57 27206
rect -257 26930 -238 27070
rect -192 27052 57 27070
rect 23341 27105 23711 27206
rect 23341 27059 23592 27105
rect 23638 27059 23711 27105
rect 23341 27052 23711 27059
rect -192 26948 -173 27052
rect 23519 26948 23711 27052
rect -192 26930 57 26948
rect -257 26794 57 26930
rect 23341 26941 23711 26948
rect 23341 26895 23592 26941
rect 23638 26895 23711 26941
rect 23341 26794 23711 26895
rect -257 25270 57 25406
rect -257 25130 -238 25270
rect -192 25252 57 25270
rect 23341 25305 23711 25406
rect 23341 25259 23592 25305
rect 23638 25259 23711 25305
rect 23341 25252 23711 25259
rect -192 25148 -173 25252
rect 23519 25148 23711 25252
rect -192 25130 57 25148
rect -257 24994 57 25130
rect 23341 25141 23711 25148
rect 23341 25095 23592 25141
rect 23638 25095 23711 25141
rect 23341 24994 23711 25095
rect -257 23470 57 23606
rect -257 23330 -238 23470
rect -192 23452 57 23470
rect 23341 23505 23711 23606
rect 23341 23459 23592 23505
rect 23638 23459 23711 23505
rect 23341 23452 23711 23459
rect -192 23348 -173 23452
rect 23519 23348 23711 23452
rect -192 23330 57 23348
rect -257 23194 57 23330
rect 23341 23341 23711 23348
rect 23341 23295 23592 23341
rect 23638 23295 23711 23341
rect 23341 23194 23711 23295
rect -257 21670 57 21806
rect -257 21530 -238 21670
rect -192 21652 57 21670
rect 23341 21705 23711 21806
rect 23341 21659 23592 21705
rect 23638 21659 23711 21705
rect 23341 21652 23711 21659
rect -192 21548 -173 21652
rect 23519 21548 23711 21652
rect -192 21530 57 21548
rect -257 21394 57 21530
rect 23341 21541 23711 21548
rect 23341 21495 23592 21541
rect 23638 21495 23711 21541
rect 23341 21394 23711 21495
rect -257 19870 57 20006
rect -257 19730 -238 19870
rect -192 19852 57 19870
rect 23341 19905 23711 20006
rect 23341 19859 23592 19905
rect 23638 19859 23711 19905
rect 23341 19852 23711 19859
rect -192 19748 -173 19852
rect 23519 19748 23711 19852
rect -192 19730 57 19748
rect -257 19594 57 19730
rect 23341 19741 23711 19748
rect 23341 19695 23592 19741
rect 23638 19695 23711 19741
rect 23341 19594 23711 19695
rect -257 18070 57 18206
rect -257 17930 -238 18070
rect -192 18052 57 18070
rect 23341 18105 23711 18206
rect 23341 18059 23592 18105
rect 23638 18059 23711 18105
rect 23341 18052 23711 18059
rect -192 17948 -173 18052
rect 23519 17948 23711 18052
rect -192 17930 57 17948
rect -257 17794 57 17930
rect 23341 17941 23711 17948
rect 23341 17895 23592 17941
rect 23638 17895 23711 17941
rect 23341 17794 23711 17895
rect -257 16270 57 16406
rect -257 16130 -238 16270
rect -192 16252 57 16270
rect 23341 16305 23711 16406
rect 23341 16259 23592 16305
rect 23638 16259 23711 16305
rect 23341 16252 23711 16259
rect -192 16148 -173 16252
rect 23519 16148 23711 16252
rect -192 16130 57 16148
rect -257 15994 57 16130
rect 23341 16141 23711 16148
rect 23341 16095 23592 16141
rect 23638 16095 23711 16141
rect 23341 15994 23711 16095
rect -257 14470 57 14606
rect -257 14330 -238 14470
rect -192 14452 57 14470
rect 23341 14505 23711 14606
rect 23341 14459 23592 14505
rect 23638 14459 23711 14505
rect 23341 14452 23711 14459
rect -192 14348 -173 14452
rect 23519 14348 23711 14452
rect -192 14330 57 14348
rect -257 14194 57 14330
rect 23341 14341 23711 14348
rect 23341 14295 23592 14341
rect 23638 14295 23711 14341
rect 23341 14194 23711 14295
rect -257 12670 57 12806
rect -257 12530 -238 12670
rect -192 12652 57 12670
rect 23341 12705 23711 12806
rect 23341 12659 23592 12705
rect 23638 12659 23711 12705
rect 23341 12652 23711 12659
rect -192 12548 -173 12652
rect 23519 12548 23711 12652
rect -192 12530 57 12548
rect -257 12394 57 12530
rect 23341 12541 23711 12548
rect 23341 12495 23592 12541
rect 23638 12495 23711 12541
rect 23341 12394 23711 12495
rect -257 10870 57 11006
rect -257 10730 -238 10870
rect -192 10852 57 10870
rect 23341 10905 23711 11006
rect 23341 10859 23592 10905
rect 23638 10859 23711 10905
rect 23341 10852 23711 10859
rect -192 10748 -173 10852
rect 23519 10748 23711 10852
rect -192 10730 57 10748
rect -257 10594 57 10730
rect 23341 10741 23711 10748
rect 23341 10695 23592 10741
rect 23638 10695 23711 10741
rect 23341 10594 23711 10695
rect -257 9070 57 9206
rect -257 8930 -238 9070
rect -192 9052 57 9070
rect 23341 9105 23711 9206
rect 23341 9059 23592 9105
rect 23638 9059 23711 9105
rect 23341 9052 23711 9059
rect -192 8948 -173 9052
rect 23519 8948 23711 9052
rect -192 8930 57 8948
rect -257 8794 57 8930
rect 23341 8941 23711 8948
rect 23341 8895 23592 8941
rect 23638 8895 23711 8941
rect 23341 8794 23711 8895
rect -257 7270 57 7406
rect -257 7130 -238 7270
rect -192 7252 57 7270
rect 23341 7305 23711 7406
rect 23341 7259 23592 7305
rect 23638 7259 23711 7305
rect 23341 7252 23711 7259
rect -192 7148 -173 7252
rect 23519 7148 23711 7252
rect -192 7130 57 7148
rect -257 6994 57 7130
rect 23341 7141 23711 7148
rect 23341 7095 23592 7141
rect 23638 7095 23711 7141
rect 23341 6994 23711 7095
rect -257 5470 57 5606
rect -257 5330 -238 5470
rect -192 5452 57 5470
rect 23341 5505 23711 5606
rect 23341 5459 23592 5505
rect 23638 5459 23711 5505
rect 23341 5452 23711 5459
rect -192 5348 -173 5452
rect 23519 5348 23711 5452
rect -192 5330 57 5348
rect -257 5194 57 5330
rect 23341 5341 23711 5348
rect 23341 5295 23592 5341
rect 23638 5295 23711 5341
rect 23341 5194 23711 5295
rect -257 3670 57 3806
rect -257 3530 -238 3670
rect -192 3652 57 3670
rect 23341 3705 23711 3806
rect 23341 3659 23592 3705
rect 23638 3659 23711 3705
rect 23341 3652 23711 3659
rect -192 3548 -173 3652
rect 23519 3548 23711 3652
rect -192 3530 57 3548
rect -257 3394 57 3530
rect 23341 3541 23711 3548
rect 23341 3495 23592 3541
rect 23638 3495 23711 3541
rect 23341 3394 23711 3495
rect -257 1870 57 2006
rect -257 1730 -238 1870
rect -192 1852 57 1870
rect 23341 1905 23711 2006
rect 23341 1859 23592 1905
rect 23638 1859 23711 1905
rect 23341 1852 23711 1859
rect -192 1748 -173 1852
rect 23519 1748 23711 1852
rect -192 1730 57 1748
rect -257 1594 57 1730
rect 23341 1741 23711 1748
rect 23341 1695 23592 1741
rect 23638 1695 23711 1741
rect 23341 1594 23711 1695
rect 23519 345 23711 391
rect 23519 299 23592 345
rect 23638 299 23711 345
rect -257 211 -173 230
rect -257 71 -238 211
rect -192 206 -173 211
rect 23519 206 23711 299
rect -192 71 57 206
rect -257 52 57 71
rect 23395 181 23711 206
rect 23395 135 23592 181
rect 23638 135 23711 181
rect 23395 52 23711 135
rect 22957 -15781 23034 -15739
rect 23181 -15781 23258 -15739
rect 22936 -15798 23056 -15781
rect 23160 -15798 23280 -15781
rect 22936 -15814 23280 -15798
rect 22936 -15860 23569 -15814
rect 22936 -15906 23291 -15860
rect 23337 -15906 23449 -15860
rect 23495 -15906 23569 -15860
rect 22936 -15952 23569 -15906
rect 22936 -15961 23280 -15952
rect 22936 -16022 23056 -15961
rect 23160 -16022 23280 -15961
rect 22936 -16401 23056 -16319
rect 23160 -16401 23280 -16319
rect 22940 -19466 23060 -19404
rect 23164 -19466 23284 -19404
rect 22940 -19475 23284 -19466
rect 22633 -19521 23284 -19475
rect 22633 -19567 22707 -19521
rect 22753 -19567 22865 -19521
rect 22911 -19567 23284 -19521
rect 22633 -19613 23284 -19567
rect 22940 -19624 23284 -19613
rect 22940 -19640 23060 -19624
rect 23164 -19640 23284 -19624
rect 22961 -19683 23038 -19640
rect 23185 -19683 23262 -19640
<< polycontact >>
rect -238 59189 -192 59329
rect 23592 59219 23638 59265
rect 23592 59055 23638 59101
rect -238 57530 -192 57670
rect 23592 57659 23638 57705
rect 23592 57495 23638 57541
rect -238 55730 -192 55870
rect 23592 55859 23638 55905
rect 23592 55695 23638 55741
rect -238 53930 -192 54070
rect 23592 54059 23638 54105
rect 23592 53895 23638 53941
rect -238 52130 -192 52270
rect 23592 52259 23638 52305
rect 23592 52095 23638 52141
rect -238 50330 -192 50470
rect 23592 50459 23638 50505
rect 23592 50295 23638 50341
rect -238 48530 -192 48670
rect 23592 48659 23638 48705
rect 23592 48495 23638 48541
rect -238 46730 -192 46870
rect 23592 46859 23638 46905
rect 23592 46695 23638 46741
rect -238 44930 -192 45070
rect 23592 45059 23638 45105
rect 23592 44895 23638 44941
rect -238 43130 -192 43270
rect 23592 43259 23638 43305
rect 23592 43095 23638 43141
rect -238 41330 -192 41470
rect 23592 41459 23638 41505
rect 23592 41295 23638 41341
rect -238 39530 -192 39670
rect 23592 39659 23638 39705
rect 23592 39495 23638 39541
rect -238 37730 -192 37870
rect 23592 37859 23638 37905
rect 23592 37695 23638 37741
rect -238 35930 -192 36070
rect 23592 36059 23638 36105
rect 23592 35895 23638 35941
rect -238 34130 -192 34270
rect 23592 34259 23638 34305
rect 23592 34095 23638 34141
rect -238 32330 -192 32470
rect 23592 32459 23638 32505
rect 23592 32295 23638 32341
rect -238 30530 -192 30670
rect 23592 30659 23638 30705
rect 23592 30495 23638 30541
rect -238 28730 -192 28870
rect 23592 28859 23638 28905
rect 23592 28695 23638 28741
rect -238 26930 -192 27070
rect 23592 27059 23638 27105
rect 23592 26895 23638 26941
rect -238 25130 -192 25270
rect 23592 25259 23638 25305
rect 23592 25095 23638 25141
rect -238 23330 -192 23470
rect 23592 23459 23638 23505
rect 23592 23295 23638 23341
rect -238 21530 -192 21670
rect 23592 21659 23638 21705
rect 23592 21495 23638 21541
rect -238 19730 -192 19870
rect 23592 19859 23638 19905
rect 23592 19695 23638 19741
rect -238 17930 -192 18070
rect 23592 18059 23638 18105
rect 23592 17895 23638 17941
rect -238 16130 -192 16270
rect 23592 16259 23638 16305
rect 23592 16095 23638 16141
rect -238 14330 -192 14470
rect 23592 14459 23638 14505
rect 23592 14295 23638 14341
rect -238 12530 -192 12670
rect 23592 12659 23638 12705
rect 23592 12495 23638 12541
rect -238 10730 -192 10870
rect 23592 10859 23638 10905
rect 23592 10695 23638 10741
rect -238 8930 -192 9070
rect 23592 9059 23638 9105
rect 23592 8895 23638 8941
rect -238 7130 -192 7270
rect 23592 7259 23638 7305
rect 23592 7095 23638 7141
rect -238 5330 -192 5470
rect 23592 5459 23638 5505
rect 23592 5295 23638 5341
rect -238 3530 -192 3670
rect 23592 3659 23638 3705
rect 23592 3495 23638 3541
rect -238 1730 -192 1870
rect 23592 1859 23638 1905
rect 23592 1695 23638 1741
rect 23592 299 23638 345
rect -238 71 -192 211
rect 23592 135 23638 181
rect 23291 -15906 23337 -15860
rect 23449 -15906 23495 -15860
rect 22707 -19567 22753 -19521
rect 22865 -19567 22911 -19521
<< metal1 >>
rect -253 59329 -177 59340
rect -253 59328 -238 59329
rect -192 59328 -177 59329
rect -253 59068 -241 59328
rect -189 59068 -177 59328
rect -253 59056 -177 59068
rect 23551 59270 23675 59310
rect 23551 59218 23587 59270
rect 23639 59218 23675 59270
rect 23551 59101 23675 59218
rect 23551 59055 23592 59101
rect 23638 59055 23675 59101
rect 23551 59052 23675 59055
rect 23551 59000 23587 59052
rect 23639 59000 23675 59052
rect 23551 58960 23675 59000
rect -253 57729 -177 57741
rect -253 57469 -241 57729
rect -189 57469 -177 57729
rect -253 57457 -177 57469
rect 23551 57733 23675 57773
rect 23551 57681 23587 57733
rect 23639 57681 23675 57733
rect 23551 57659 23592 57681
rect 23638 57659 23675 57681
rect 23551 57541 23675 57659
rect 23551 57515 23592 57541
rect 23638 57515 23675 57541
rect 23551 57463 23587 57515
rect 23639 57463 23675 57515
rect 23551 57423 23675 57463
rect -253 55930 -177 55942
rect -253 55670 -241 55930
rect -189 55670 -177 55930
rect -253 55658 -177 55670
rect 23551 55933 23675 55973
rect 23551 55881 23587 55933
rect 23639 55881 23675 55933
rect 23551 55859 23592 55881
rect 23638 55859 23675 55881
rect 23551 55741 23675 55859
rect 23551 55715 23592 55741
rect 23638 55715 23675 55741
rect 23551 55663 23587 55715
rect 23639 55663 23675 55715
rect 23551 55623 23675 55663
rect -253 54130 -177 54142
rect -253 53870 -241 54130
rect -189 53870 -177 54130
rect -253 53858 -177 53870
rect 23551 54133 23675 54173
rect 23551 54081 23587 54133
rect 23639 54081 23675 54133
rect 23551 54059 23592 54081
rect 23638 54059 23675 54081
rect 23551 53941 23675 54059
rect 23551 53915 23592 53941
rect 23638 53915 23675 53941
rect 23551 53863 23587 53915
rect 23639 53863 23675 53915
rect 23551 53823 23675 53863
rect -253 52330 -177 52342
rect -253 52070 -241 52330
rect -189 52070 -177 52330
rect -253 52058 -177 52070
rect 23551 52333 23675 52373
rect 23551 52281 23587 52333
rect 23639 52281 23675 52333
rect 23551 52259 23592 52281
rect 23638 52259 23675 52281
rect 23551 52141 23675 52259
rect 23551 52115 23592 52141
rect 23638 52115 23675 52141
rect 23551 52063 23587 52115
rect 23639 52063 23675 52115
rect 23551 52023 23675 52063
rect -253 50529 -177 50541
rect -253 50269 -241 50529
rect -189 50269 -177 50529
rect -253 50257 -177 50269
rect 23551 50533 23675 50573
rect 23551 50481 23587 50533
rect 23639 50500 23675 50533
rect 23639 50481 24098 50500
rect 23551 50459 23592 50481
rect 23638 50459 24098 50481
rect 23551 50341 24098 50459
rect 23551 50315 23592 50341
rect 23638 50315 24098 50341
rect 23551 50263 23587 50315
rect 23639 50300 24098 50315
rect 23639 50263 23675 50300
rect 23551 50223 23675 50263
rect -253 48730 -177 48742
rect -253 48470 -241 48730
rect -189 48470 -177 48730
rect -253 48458 -177 48470
rect 23551 48733 23675 48773
rect 23551 48681 23587 48733
rect 23639 48681 23675 48733
rect 23551 48659 23592 48681
rect 23638 48659 23675 48681
rect 23551 48541 23675 48659
rect 23551 48515 23592 48541
rect 23638 48515 23675 48541
rect 23551 48463 23587 48515
rect 23639 48463 23675 48515
rect 23551 48423 23675 48463
rect -253 46931 -177 46943
rect -253 46671 -241 46931
rect -189 46671 -177 46931
rect -253 46659 -177 46671
rect 23551 46933 23675 46973
rect 23551 46881 23587 46933
rect 23639 46881 23675 46933
rect 23551 46859 23592 46881
rect 23638 46859 23675 46881
rect 23551 46741 23675 46859
rect 23551 46715 23592 46741
rect 23638 46715 23675 46741
rect 23551 46663 23587 46715
rect 23639 46663 23675 46715
rect 23551 46623 23675 46663
rect -253 45130 -177 45142
rect -253 44870 -241 45130
rect -189 44870 -177 45130
rect -253 44858 -177 44870
rect 23551 45133 23675 45173
rect 23551 45081 23587 45133
rect 23639 45081 23675 45133
rect 23551 45059 23592 45081
rect 23638 45059 23675 45081
rect 23551 44941 23675 45059
rect 23551 44915 23592 44941
rect 23638 44915 23675 44941
rect 23551 44863 23587 44915
rect 23639 44863 23675 44915
rect 23551 44823 23675 44863
rect -253 43330 -177 43342
rect -253 43070 -241 43330
rect -189 43070 -177 43330
rect -253 43058 -177 43070
rect 23551 43333 23675 43373
rect 23551 43281 23587 43333
rect 23639 43281 23675 43333
rect 23551 43259 23592 43281
rect 23638 43259 23675 43281
rect 23551 43141 23675 43259
rect 23551 43115 23592 43141
rect 23638 43115 23675 43141
rect 23551 43063 23587 43115
rect 23639 43063 23675 43115
rect 23551 43023 23675 43063
rect -253 41530 -177 41542
rect -253 41270 -241 41530
rect -189 41270 -177 41530
rect -253 41258 -177 41270
rect 23551 41533 23675 41573
rect 23551 41481 23587 41533
rect 23639 41481 23675 41533
rect 23551 41459 23592 41481
rect 23638 41459 23675 41481
rect 23551 41341 23675 41459
rect 23551 41315 23592 41341
rect 23638 41315 23675 41341
rect 23551 41263 23587 41315
rect 23639 41263 23675 41315
rect 23551 41223 23675 41263
rect -253 39730 -177 39742
rect -253 39470 -241 39730
rect -189 39470 -177 39730
rect -253 39458 -177 39470
rect 23551 39733 23675 39773
rect 23551 39681 23587 39733
rect 23639 39681 23675 39733
rect 23551 39659 23592 39681
rect 23638 39659 23675 39681
rect 23551 39541 23675 39659
rect 23551 39515 23592 39541
rect 23638 39515 23675 39541
rect 23551 39463 23587 39515
rect 23639 39463 23675 39515
rect 23551 39423 23675 39463
rect -253 37930 -177 37942
rect -253 37670 -241 37930
rect -189 37670 -177 37930
rect -253 37658 -177 37670
rect 23551 37933 23675 37973
rect 23551 37881 23587 37933
rect 23639 37881 23675 37933
rect 23551 37859 23592 37881
rect 23638 37859 23675 37881
rect 23551 37741 23675 37859
rect 23551 37715 23592 37741
rect 23638 37715 23675 37741
rect 23551 37663 23587 37715
rect 23639 37663 23675 37715
rect 23551 37623 23675 37663
rect -253 36130 -177 36142
rect -253 35870 -241 36130
rect -189 35870 -177 36130
rect -253 35858 -177 35870
rect 23551 36133 23675 36173
rect 23551 36081 23587 36133
rect 23639 36081 23675 36133
rect 23551 36059 23592 36081
rect 23638 36059 23675 36081
rect 23551 35941 23675 36059
rect 23551 35915 23592 35941
rect 23638 35915 23675 35941
rect 23551 35863 23587 35915
rect 23639 35863 23675 35915
rect 23551 35823 23675 35863
rect -253 34330 -177 34342
rect -253 34070 -241 34330
rect -189 34070 -177 34330
rect -253 34058 -177 34070
rect 23551 34333 23675 34373
rect 23551 34281 23587 34333
rect 23639 34281 23675 34333
rect 23551 34259 23592 34281
rect 23638 34259 23675 34281
rect 23551 34141 23675 34259
rect 23551 34115 23592 34141
rect 23638 34115 23675 34141
rect 23551 34063 23587 34115
rect 23639 34063 23675 34115
rect 23551 34023 23675 34063
rect -253 32530 -177 32542
rect -253 32270 -241 32530
rect -189 32270 -177 32530
rect -253 32258 -177 32270
rect 23551 32533 23675 32573
rect 23551 32481 23587 32533
rect 23639 32481 23675 32533
rect 23551 32459 23592 32481
rect 23638 32459 23675 32481
rect 23551 32341 23675 32459
rect 23551 32315 23592 32341
rect 23638 32315 23675 32341
rect 23551 32263 23587 32315
rect 23639 32263 23675 32315
rect 23551 32223 23675 32263
rect -253 30730 -177 30742
rect -253 30470 -241 30730
rect -189 30470 -177 30730
rect -253 30458 -177 30470
rect 23551 30733 23675 30773
rect 23551 30681 23587 30733
rect 23639 30681 23675 30733
rect 23551 30659 23592 30681
rect 23638 30659 23675 30681
rect 23551 30541 23675 30659
rect 23551 30515 23592 30541
rect 23638 30515 23675 30541
rect 23551 30463 23587 30515
rect 23639 30463 23675 30515
rect 23551 30423 23675 30463
rect -253 28930 -177 28942
rect -253 28670 -241 28930
rect -189 28670 -177 28930
rect -253 28658 -177 28670
rect 23551 28933 23675 28973
rect 23551 28881 23587 28933
rect 23639 28881 23675 28933
rect 23551 28859 23592 28881
rect 23638 28859 23675 28881
rect 23551 28741 23675 28859
rect 23551 28715 23592 28741
rect 23638 28715 23675 28741
rect 23551 28663 23587 28715
rect 23639 28663 23675 28715
rect 23551 28623 23675 28663
rect -253 27130 -177 27142
rect -253 26870 -241 27130
rect -189 26870 -177 27130
rect -253 26858 -177 26870
rect 23551 27133 23675 27173
rect 23551 27081 23587 27133
rect 23639 27081 23675 27133
rect 23551 27059 23592 27081
rect 23638 27059 23675 27081
rect 23551 26941 23675 27059
rect 23551 26915 23592 26941
rect 23638 26915 23675 26941
rect 23551 26863 23587 26915
rect 23639 26863 23675 26915
rect 23551 26823 23675 26863
rect -253 25330 -177 25342
rect -253 25070 -241 25330
rect -189 25070 -177 25330
rect -253 25058 -177 25070
rect 23551 25337 23675 25377
rect 23551 25285 23587 25337
rect 23639 25285 23675 25337
rect 23551 25259 23592 25285
rect 23638 25259 23675 25285
rect 23551 25141 23675 25259
rect 23551 25119 23592 25141
rect 23638 25119 23675 25141
rect 23551 25067 23587 25119
rect 23639 25067 23675 25119
rect 23551 25027 23675 25067
rect -257 23530 -181 23542
rect -257 23270 -245 23530
rect -193 23470 -181 23530
rect -192 23330 -181 23470
rect -193 23270 -181 23330
rect -257 23258 -181 23270
rect 23551 23533 23675 23573
rect 23551 23481 23587 23533
rect 23639 23481 23675 23533
rect 23551 23459 23592 23481
rect 23638 23459 23675 23481
rect 23551 23341 23675 23459
rect 23551 23315 23592 23341
rect 23638 23315 23675 23341
rect 23551 23263 23587 23315
rect 23639 23263 23675 23315
rect 23551 23223 23675 23263
rect -253 21730 -177 21742
rect -253 21470 -241 21730
rect -189 21470 -177 21730
rect -253 21458 -177 21470
rect 23551 21737 23675 21777
rect 23551 21685 23587 21737
rect 23639 21685 23675 21737
rect 23551 21659 23592 21685
rect 23638 21659 23675 21685
rect 23551 21541 23675 21659
rect 23551 21519 23592 21541
rect 23638 21519 23675 21541
rect 23551 21467 23587 21519
rect 23639 21467 23675 21519
rect 23551 21427 23675 21467
rect -253 19930 -177 19942
rect -253 19670 -241 19930
rect -189 19670 -177 19930
rect -253 19658 -177 19670
rect 23551 19933 23675 19973
rect 23551 19881 23587 19933
rect 23639 19881 23675 19933
rect 23551 19859 23592 19881
rect 23638 19859 23675 19881
rect 23551 19741 23675 19859
rect 23551 19715 23592 19741
rect 23638 19715 23675 19741
rect 23551 19663 23587 19715
rect 23639 19663 23675 19715
rect 23551 19623 23675 19663
rect -253 18130 -177 18142
rect -253 17870 -241 18130
rect -189 17870 -177 18130
rect -253 17858 -177 17870
rect 23551 18137 23675 18177
rect 23551 18085 23587 18137
rect 23639 18085 23675 18137
rect 23551 18059 23592 18085
rect 23638 18059 23675 18085
rect 23551 17941 23675 18059
rect 23551 17919 23592 17941
rect 23638 17919 23675 17941
rect 23551 17867 23587 17919
rect 23639 17867 23675 17919
rect 23551 17827 23675 17867
rect -253 16330 -177 16342
rect -253 16070 -241 16330
rect -189 16070 -177 16330
rect -253 16058 -177 16070
rect 23551 16333 23675 16373
rect 23551 16281 23587 16333
rect 23639 16281 23675 16333
rect 23551 16259 23592 16281
rect 23638 16259 23675 16281
rect 23551 16141 23675 16259
rect 23551 16115 23592 16141
rect 23638 16115 23675 16141
rect 23551 16063 23587 16115
rect 23639 16063 23675 16115
rect 23551 16023 23675 16063
rect -253 14530 -177 14542
rect -253 14270 -241 14530
rect -189 14270 -177 14530
rect -253 14258 -177 14270
rect 23551 14537 23675 14577
rect 23551 14485 23587 14537
rect 23639 14485 23675 14537
rect 23551 14459 23592 14485
rect 23638 14459 23675 14485
rect 23551 14341 23675 14459
rect 23551 14319 23592 14341
rect 23638 14319 23675 14341
rect 23551 14267 23587 14319
rect 23639 14267 23675 14319
rect 23551 14227 23675 14267
rect -253 12730 -177 12742
rect -253 12470 -241 12730
rect -189 12470 -177 12730
rect -253 12458 -177 12470
rect 23551 12733 23675 12773
rect 23551 12681 23587 12733
rect 23639 12681 23675 12733
rect 23551 12659 23592 12681
rect 23638 12659 23675 12681
rect 23551 12541 23675 12659
rect 23551 12515 23592 12541
rect 23638 12515 23675 12541
rect 23551 12463 23587 12515
rect 23639 12463 23675 12515
rect 23551 12423 23675 12463
rect -253 10930 -177 10942
rect -253 10670 -241 10930
rect -189 10670 -177 10930
rect -253 10658 -177 10670
rect 23551 10937 23675 10977
rect 23551 10885 23587 10937
rect 23639 10885 23675 10937
rect 23551 10859 23592 10885
rect 23638 10859 23675 10885
rect 23551 10741 23675 10859
rect 23551 10719 23592 10741
rect 23638 10719 23675 10741
rect 23551 10667 23587 10719
rect 23639 10667 23675 10719
rect 23551 10627 23675 10667
rect -253 9130 -177 9142
rect -253 8870 -241 9130
rect -189 8870 -177 9130
rect -253 8858 -177 8870
rect 23551 9133 23675 9173
rect 23551 9081 23587 9133
rect 23639 9081 23675 9133
rect 23551 9059 23592 9081
rect 23638 9059 23675 9081
rect 23551 8941 23675 9059
rect 23551 8915 23592 8941
rect 23638 8915 23675 8941
rect 23551 8863 23587 8915
rect 23639 8863 23675 8915
rect 23551 8823 23675 8863
rect -253 7330 -177 7342
rect -253 7070 -241 7330
rect -189 7070 -177 7330
rect -253 7058 -177 7070
rect 23551 7337 23675 7377
rect 23551 7285 23587 7337
rect 23639 7285 23675 7337
rect 23551 7259 23592 7285
rect 23638 7259 23675 7285
rect 23551 7141 23675 7259
rect 23551 7119 23592 7141
rect 23638 7119 23675 7141
rect 23551 7067 23587 7119
rect 23639 7067 23675 7119
rect 23551 7027 23675 7067
rect -253 5530 -177 5542
rect -253 5270 -241 5530
rect -189 5270 -177 5530
rect -253 5258 -177 5270
rect 23551 5533 23675 5573
rect 23551 5481 23587 5533
rect 23639 5481 23675 5533
rect 23551 5459 23592 5481
rect 23638 5459 23675 5481
rect 23551 5341 23675 5459
rect 23551 5315 23592 5341
rect 23638 5315 23675 5341
rect 23551 5263 23587 5315
rect 23639 5263 23675 5315
rect 23551 5223 23675 5263
rect -253 3730 -177 3742
rect -253 3470 -241 3730
rect -189 3470 -177 3730
rect -253 3458 -177 3470
rect 23551 3737 23675 3777
rect 23551 3685 23587 3737
rect 23639 3685 23675 3737
rect 23551 3659 23592 3685
rect 23638 3659 23675 3685
rect 23551 3541 23675 3659
rect 23551 3519 23592 3541
rect 23638 3519 23675 3541
rect 23551 3467 23587 3519
rect 23639 3467 23675 3519
rect 23551 3427 23675 3467
rect -253 1930 -177 1942
rect -253 1670 -241 1930
rect -189 1670 -177 1930
rect -253 1658 -177 1670
rect 23551 1933 23675 1973
rect 23551 1881 23587 1933
rect 23639 1881 23675 1933
rect 23551 1859 23592 1881
rect 23638 1859 23675 1881
rect 23551 1741 23675 1859
rect 23551 1715 23592 1741
rect 23638 1715 23675 1741
rect 23551 1663 23587 1715
rect 23639 1663 23675 1715
rect 23551 1623 23675 1663
rect 23551 400 23675 440
rect 23551 348 23587 400
rect 23639 348 23675 400
rect 23551 345 23675 348
rect 23551 299 23592 345
rect 23638 299 23675 345
rect -255 211 -179 280
rect -255 71 -238 211
rect -192 71 -179 211
rect 23551 182 23675 299
rect 23551 130 23587 182
rect 23639 130 23675 182
rect 23551 90 23675 130
rect -255 -317 -179 71
rect -255 -487 66 -317
rect 22970 -6200 23184 -4838
rect 22472 -11894 23031 -11774
rect 22472 -13621 22588 -11894
rect 23211 -12293 23453 -11996
rect 22472 -13741 23603 -13621
rect 22834 -14599 23266 -14562
rect 22834 -14645 22869 -14599
rect 22915 -14645 23027 -14599
rect 23073 -14645 23185 -14599
rect 23231 -14645 23266 -14599
rect 22834 -14682 23266 -14645
rect 23049 -15809 23166 -15424
rect 22648 -15884 23166 -15809
rect 23486 -15823 23603 -13741
rect 22648 -19484 22720 -15884
rect 23049 -16147 23166 -15884
rect 23256 -15860 23603 -15823
rect 23256 -15906 23291 -15860
rect 23337 -15906 23449 -15860
rect 23495 -15906 23603 -15860
rect 23256 -15943 23603 -15906
rect 22825 -16543 22942 -16269
rect 23273 -16543 23390 -16269
rect 22825 -16594 23390 -16543
rect 22825 -16640 22926 -16594
rect 22972 -16640 23084 -16594
rect 23130 -16640 23242 -16594
rect 23288 -16640 23390 -16594
rect 22825 -16691 23390 -16640
rect 22825 -18488 22942 -16691
rect 22648 -19521 22946 -19484
rect 22648 -19567 22707 -19521
rect 22753 -19567 22865 -19521
rect 22911 -19567 22946 -19521
rect 22648 -19604 22946 -19567
rect 23054 -19830 23170 -18443
rect 23273 -18488 23390 -16691
rect 22830 -22882 22946 -21688
rect 23278 -22882 23394 -21688
rect 22717 -22919 22946 -22882
rect 22717 -22965 22751 -22919
rect 22797 -22965 22946 -22919
rect 22717 -23002 22946 -22965
rect 23049 -23165 23179 -22898
rect 23261 -22919 23394 -22882
rect 23261 -22965 23295 -22919
rect 23341 -22965 23394 -22919
rect 23261 -23002 23394 -22965
rect 23001 -25410 23223 -23165
<< via1 >>
rect -241 59189 -238 59328
rect -238 59189 -192 59328
rect -192 59189 -189 59328
rect -241 59068 -189 59189
rect 23587 59265 23639 59270
rect 23587 59219 23592 59265
rect 23592 59219 23638 59265
rect 23638 59219 23639 59265
rect 23587 59218 23639 59219
rect 23587 59000 23639 59052
rect -241 57670 -189 57729
rect -241 57530 -238 57670
rect -238 57530 -192 57670
rect -192 57530 -189 57670
rect -241 57469 -189 57530
rect 23587 57705 23639 57733
rect 23587 57681 23592 57705
rect 23592 57681 23638 57705
rect 23638 57681 23639 57705
rect 23587 57495 23592 57515
rect 23592 57495 23638 57515
rect 23638 57495 23639 57515
rect 23587 57463 23639 57495
rect -241 55870 -189 55930
rect -241 55730 -238 55870
rect -238 55730 -192 55870
rect -192 55730 -189 55870
rect -241 55670 -189 55730
rect 23587 55905 23639 55933
rect 23587 55881 23592 55905
rect 23592 55881 23638 55905
rect 23638 55881 23639 55905
rect 23587 55695 23592 55715
rect 23592 55695 23638 55715
rect 23638 55695 23639 55715
rect 23587 55663 23639 55695
rect -241 54070 -189 54130
rect -241 53930 -238 54070
rect -238 53930 -192 54070
rect -192 53930 -189 54070
rect -241 53870 -189 53930
rect 23587 54105 23639 54133
rect 23587 54081 23592 54105
rect 23592 54081 23638 54105
rect 23638 54081 23639 54105
rect 23587 53895 23592 53915
rect 23592 53895 23638 53915
rect 23638 53895 23639 53915
rect 23587 53863 23639 53895
rect -241 52270 -189 52330
rect -241 52130 -238 52270
rect -238 52130 -192 52270
rect -192 52130 -189 52270
rect -241 52070 -189 52130
rect 23587 52305 23639 52333
rect 23587 52281 23592 52305
rect 23592 52281 23638 52305
rect 23638 52281 23639 52305
rect 23587 52095 23592 52115
rect 23592 52095 23638 52115
rect 23638 52095 23639 52115
rect 23587 52063 23639 52095
rect -241 50470 -189 50529
rect -241 50330 -238 50470
rect -238 50330 -192 50470
rect -192 50330 -189 50470
rect -241 50269 -189 50330
rect 23587 50505 23639 50533
rect 23587 50481 23592 50505
rect 23592 50481 23638 50505
rect 23638 50481 23639 50505
rect 23587 50295 23592 50315
rect 23592 50295 23638 50315
rect 23638 50295 23639 50315
rect 23587 50263 23639 50295
rect -241 48670 -189 48730
rect -241 48530 -238 48670
rect -238 48530 -192 48670
rect -192 48530 -189 48670
rect -241 48470 -189 48530
rect 23587 48705 23639 48733
rect 23587 48681 23592 48705
rect 23592 48681 23638 48705
rect 23638 48681 23639 48705
rect 23587 48495 23592 48515
rect 23592 48495 23638 48515
rect 23638 48495 23639 48515
rect 23587 48463 23639 48495
rect -241 46870 -189 46931
rect -241 46730 -238 46870
rect -238 46730 -192 46870
rect -192 46730 -189 46870
rect -241 46671 -189 46730
rect 23587 46905 23639 46933
rect 23587 46881 23592 46905
rect 23592 46881 23638 46905
rect 23638 46881 23639 46905
rect 23587 46695 23592 46715
rect 23592 46695 23638 46715
rect 23638 46695 23639 46715
rect 23587 46663 23639 46695
rect -241 45070 -189 45130
rect -241 44930 -238 45070
rect -238 44930 -192 45070
rect -192 44930 -189 45070
rect -241 44870 -189 44930
rect 23587 45105 23639 45133
rect 23587 45081 23592 45105
rect 23592 45081 23638 45105
rect 23638 45081 23639 45105
rect 23587 44895 23592 44915
rect 23592 44895 23638 44915
rect 23638 44895 23639 44915
rect 23587 44863 23639 44895
rect -241 43270 -189 43330
rect -241 43130 -238 43270
rect -238 43130 -192 43270
rect -192 43130 -189 43270
rect -241 43070 -189 43130
rect 23587 43305 23639 43333
rect 23587 43281 23592 43305
rect 23592 43281 23638 43305
rect 23638 43281 23639 43305
rect 23587 43095 23592 43115
rect 23592 43095 23638 43115
rect 23638 43095 23639 43115
rect 23587 43063 23639 43095
rect -241 41470 -189 41530
rect -241 41330 -238 41470
rect -238 41330 -192 41470
rect -192 41330 -189 41470
rect -241 41270 -189 41330
rect 23587 41505 23639 41533
rect 23587 41481 23592 41505
rect 23592 41481 23638 41505
rect 23638 41481 23639 41505
rect 23587 41295 23592 41315
rect 23592 41295 23638 41315
rect 23638 41295 23639 41315
rect 23587 41263 23639 41295
rect -241 39670 -189 39730
rect -241 39530 -238 39670
rect -238 39530 -192 39670
rect -192 39530 -189 39670
rect -241 39470 -189 39530
rect 23587 39705 23639 39733
rect 23587 39681 23592 39705
rect 23592 39681 23638 39705
rect 23638 39681 23639 39705
rect 23587 39495 23592 39515
rect 23592 39495 23638 39515
rect 23638 39495 23639 39515
rect 23587 39463 23639 39495
rect -241 37870 -189 37930
rect -241 37730 -238 37870
rect -238 37730 -192 37870
rect -192 37730 -189 37870
rect -241 37670 -189 37730
rect 23587 37905 23639 37933
rect 23587 37881 23592 37905
rect 23592 37881 23638 37905
rect 23638 37881 23639 37905
rect 23587 37695 23592 37715
rect 23592 37695 23638 37715
rect 23638 37695 23639 37715
rect 23587 37663 23639 37695
rect -241 36070 -189 36130
rect -241 35930 -238 36070
rect -238 35930 -192 36070
rect -192 35930 -189 36070
rect -241 35870 -189 35930
rect 23587 36105 23639 36133
rect 23587 36081 23592 36105
rect 23592 36081 23638 36105
rect 23638 36081 23639 36105
rect 23587 35895 23592 35915
rect 23592 35895 23638 35915
rect 23638 35895 23639 35915
rect 23587 35863 23639 35895
rect -241 34270 -189 34330
rect -241 34130 -238 34270
rect -238 34130 -192 34270
rect -192 34130 -189 34270
rect -241 34070 -189 34130
rect 23587 34305 23639 34333
rect 23587 34281 23592 34305
rect 23592 34281 23638 34305
rect 23638 34281 23639 34305
rect 23587 34095 23592 34115
rect 23592 34095 23638 34115
rect 23638 34095 23639 34115
rect 23587 34063 23639 34095
rect -241 32470 -189 32530
rect -241 32330 -238 32470
rect -238 32330 -192 32470
rect -192 32330 -189 32470
rect -241 32270 -189 32330
rect 23587 32505 23639 32533
rect 23587 32481 23592 32505
rect 23592 32481 23638 32505
rect 23638 32481 23639 32505
rect 23587 32295 23592 32315
rect 23592 32295 23638 32315
rect 23638 32295 23639 32315
rect 23587 32263 23639 32295
rect -241 30670 -189 30730
rect -241 30530 -238 30670
rect -238 30530 -192 30670
rect -192 30530 -189 30670
rect -241 30470 -189 30530
rect 23587 30705 23639 30733
rect 23587 30681 23592 30705
rect 23592 30681 23638 30705
rect 23638 30681 23639 30705
rect 23587 30495 23592 30515
rect 23592 30495 23638 30515
rect 23638 30495 23639 30515
rect 23587 30463 23639 30495
rect -241 28870 -189 28930
rect -241 28730 -238 28870
rect -238 28730 -192 28870
rect -192 28730 -189 28870
rect -241 28670 -189 28730
rect 23587 28905 23639 28933
rect 23587 28881 23592 28905
rect 23592 28881 23638 28905
rect 23638 28881 23639 28905
rect 23587 28695 23592 28715
rect 23592 28695 23638 28715
rect 23638 28695 23639 28715
rect 23587 28663 23639 28695
rect -241 27070 -189 27130
rect -241 26930 -238 27070
rect -238 26930 -192 27070
rect -192 26930 -189 27070
rect -241 26870 -189 26930
rect 23587 27105 23639 27133
rect 23587 27081 23592 27105
rect 23592 27081 23638 27105
rect 23638 27081 23639 27105
rect 23587 26895 23592 26915
rect 23592 26895 23638 26915
rect 23638 26895 23639 26915
rect 23587 26863 23639 26895
rect -241 25270 -189 25330
rect -241 25130 -238 25270
rect -238 25130 -192 25270
rect -192 25130 -189 25270
rect -241 25070 -189 25130
rect 23587 25305 23639 25337
rect 23587 25285 23592 25305
rect 23592 25285 23638 25305
rect 23638 25285 23639 25305
rect 23587 25095 23592 25119
rect 23592 25095 23638 25119
rect 23638 25095 23639 25119
rect 23587 25067 23639 25095
rect -245 23470 -193 23530
rect -245 23330 -238 23470
rect -238 23330 -193 23470
rect -245 23270 -193 23330
rect 23587 23505 23639 23533
rect 23587 23481 23592 23505
rect 23592 23481 23638 23505
rect 23638 23481 23639 23505
rect 23587 23295 23592 23315
rect 23592 23295 23638 23315
rect 23638 23295 23639 23315
rect 23587 23263 23639 23295
rect -241 21670 -189 21730
rect -241 21530 -238 21670
rect -238 21530 -192 21670
rect -192 21530 -189 21670
rect -241 21470 -189 21530
rect 23587 21705 23639 21737
rect 23587 21685 23592 21705
rect 23592 21685 23638 21705
rect 23638 21685 23639 21705
rect 23587 21495 23592 21519
rect 23592 21495 23638 21519
rect 23638 21495 23639 21519
rect 23587 21467 23639 21495
rect -241 19870 -189 19930
rect -241 19730 -238 19870
rect -238 19730 -192 19870
rect -192 19730 -189 19870
rect -241 19670 -189 19730
rect 23587 19905 23639 19933
rect 23587 19881 23592 19905
rect 23592 19881 23638 19905
rect 23638 19881 23639 19905
rect 23587 19695 23592 19715
rect 23592 19695 23638 19715
rect 23638 19695 23639 19715
rect 23587 19663 23639 19695
rect -241 18070 -189 18130
rect -241 17930 -238 18070
rect -238 17930 -192 18070
rect -192 17930 -189 18070
rect -241 17870 -189 17930
rect 23587 18105 23639 18137
rect 23587 18085 23592 18105
rect 23592 18085 23638 18105
rect 23638 18085 23639 18105
rect 23587 17895 23592 17919
rect 23592 17895 23638 17919
rect 23638 17895 23639 17919
rect 23587 17867 23639 17895
rect -241 16270 -189 16330
rect -241 16130 -238 16270
rect -238 16130 -192 16270
rect -192 16130 -189 16270
rect -241 16070 -189 16130
rect 23587 16305 23639 16333
rect 23587 16281 23592 16305
rect 23592 16281 23638 16305
rect 23638 16281 23639 16305
rect 23587 16095 23592 16115
rect 23592 16095 23638 16115
rect 23638 16095 23639 16115
rect 23587 16063 23639 16095
rect -241 14470 -189 14530
rect -241 14330 -238 14470
rect -238 14330 -192 14470
rect -192 14330 -189 14470
rect -241 14270 -189 14330
rect 23587 14505 23639 14537
rect 23587 14485 23592 14505
rect 23592 14485 23638 14505
rect 23638 14485 23639 14505
rect 23587 14295 23592 14319
rect 23592 14295 23638 14319
rect 23638 14295 23639 14319
rect 23587 14267 23639 14295
rect -241 12670 -189 12730
rect -241 12530 -238 12670
rect -238 12530 -192 12670
rect -192 12530 -189 12670
rect -241 12470 -189 12530
rect 23587 12705 23639 12733
rect 23587 12681 23592 12705
rect 23592 12681 23638 12705
rect 23638 12681 23639 12705
rect 23587 12495 23592 12515
rect 23592 12495 23638 12515
rect 23638 12495 23639 12515
rect 23587 12463 23639 12495
rect -241 10870 -189 10930
rect -241 10730 -238 10870
rect -238 10730 -192 10870
rect -192 10730 -189 10870
rect -241 10670 -189 10730
rect 23587 10905 23639 10937
rect 23587 10885 23592 10905
rect 23592 10885 23638 10905
rect 23638 10885 23639 10905
rect 23587 10695 23592 10719
rect 23592 10695 23638 10719
rect 23638 10695 23639 10719
rect 23587 10667 23639 10695
rect -241 9070 -189 9130
rect -241 8930 -238 9070
rect -238 8930 -192 9070
rect -192 8930 -189 9070
rect -241 8870 -189 8930
rect 23587 9105 23639 9133
rect 23587 9081 23592 9105
rect 23592 9081 23638 9105
rect 23638 9081 23639 9105
rect 23587 8895 23592 8915
rect 23592 8895 23638 8915
rect 23638 8895 23639 8915
rect 23587 8863 23639 8895
rect -241 7270 -189 7330
rect -241 7130 -238 7270
rect -238 7130 -192 7270
rect -192 7130 -189 7270
rect -241 7070 -189 7130
rect 23587 7305 23639 7337
rect 23587 7285 23592 7305
rect 23592 7285 23638 7305
rect 23638 7285 23639 7305
rect 23587 7095 23592 7119
rect 23592 7095 23638 7119
rect 23638 7095 23639 7119
rect 23587 7067 23639 7095
rect -241 5470 -189 5530
rect -241 5330 -238 5470
rect -238 5330 -192 5470
rect -192 5330 -189 5470
rect -241 5270 -189 5330
rect 23587 5505 23639 5533
rect 23587 5481 23592 5505
rect 23592 5481 23638 5505
rect 23638 5481 23639 5505
rect 23587 5295 23592 5315
rect 23592 5295 23638 5315
rect 23638 5295 23639 5315
rect 23587 5263 23639 5295
rect -241 3670 -189 3730
rect -241 3530 -238 3670
rect -238 3530 -192 3670
rect -192 3530 -189 3670
rect -241 3470 -189 3530
rect 23587 3705 23639 3737
rect 23587 3685 23592 3705
rect 23592 3685 23638 3705
rect 23638 3685 23639 3705
rect 23587 3495 23592 3519
rect 23592 3495 23638 3519
rect 23638 3495 23639 3519
rect 23587 3467 23639 3495
rect -241 1870 -189 1930
rect -241 1730 -238 1870
rect -238 1730 -192 1870
rect -192 1730 -189 1870
rect -241 1670 -189 1730
rect 23587 1905 23639 1933
rect 23587 1881 23592 1905
rect 23592 1881 23638 1905
rect 23638 1881 23639 1905
rect 23587 1695 23592 1715
rect 23592 1695 23638 1715
rect 23638 1695 23639 1715
rect 23587 1663 23639 1695
rect 23587 348 23639 400
rect 23587 181 23639 182
rect 23587 135 23592 181
rect 23592 135 23638 181
rect 23638 135 23639 181
rect 23587 130 23639 135
<< metal2 >>
rect -253 59328 -177 59340
rect -253 59068 -241 59328
rect -189 59068 -177 59328
rect -253 57729 -177 59068
rect -253 57469 -241 57729
rect -189 57469 -177 57729
rect -253 55930 -177 57469
rect 23550 59270 23675 59310
rect 23550 59218 23587 59270
rect 23639 59218 23675 59270
rect 23550 59052 23675 59218
rect 23550 59000 23587 59052
rect 23639 59000 23675 59052
rect 23550 57733 23675 59000
rect 23550 57681 23587 57733
rect 23639 57681 23675 57733
rect 23550 57515 23675 57681
rect 23550 57463 23587 57515
rect 23639 57463 23675 57515
rect 23550 57369 23675 57463
rect -253 55670 -241 55930
rect -189 55670 -177 55930
rect -253 54130 -177 55670
rect -253 53870 -241 54130
rect -189 53870 -177 54130
rect -253 52330 -177 53870
rect -253 52070 -241 52330
rect -189 52070 -177 52330
rect -253 50529 -177 52070
rect -253 50269 -241 50529
rect -189 50269 -177 50529
rect -253 48730 -177 50269
rect -253 48470 -241 48730
rect -189 48470 -177 48730
rect -253 46931 -177 48470
rect -253 46671 -241 46931
rect -189 46671 -177 46931
rect -253 45130 -177 46671
rect -253 44870 -241 45130
rect -189 44870 -177 45130
rect -253 43330 -177 44870
rect -253 43070 -241 43330
rect -189 43070 -177 43330
rect -253 41530 -177 43070
rect -253 41270 -241 41530
rect -189 41270 -177 41530
rect -253 39730 -177 41270
rect -253 39470 -241 39730
rect -189 39470 -177 39730
rect -253 37930 -177 39470
rect -253 37670 -241 37930
rect -189 37670 -177 37930
rect -253 36130 -177 37670
rect -253 35870 -241 36130
rect -189 35870 -177 36130
rect -253 34330 -177 35870
rect -253 34070 -241 34330
rect -189 34070 -177 34330
rect -253 32530 -177 34070
rect -253 32270 -241 32530
rect -189 32270 -177 32530
rect -253 30730 -177 32270
rect -253 30470 -241 30730
rect -189 30470 -177 30730
rect -253 28930 -177 30470
rect -253 28670 -241 28930
rect -189 28670 -177 28930
rect -253 27130 -177 28670
rect -253 26870 -241 27130
rect -189 26870 -177 27130
rect -253 25330 -177 26870
rect -253 25070 -241 25330
rect -189 25070 -177 25330
rect -253 23542 -177 25070
rect -257 23530 -177 23542
rect -257 23270 -245 23530
rect -193 23270 -177 23530
rect -257 23258 -177 23270
rect -253 21730 -177 23258
rect -253 21470 -241 21730
rect -189 21470 -177 21730
rect -253 19930 -177 21470
rect -253 19670 -241 19930
rect -189 19670 -177 19930
rect -253 18130 -177 19670
rect -253 17870 -241 18130
rect -189 17870 -177 18130
rect -253 16330 -177 17870
rect -253 16070 -241 16330
rect -189 16070 -177 16330
rect -253 14530 -177 16070
rect -253 14270 -241 14530
rect -189 14270 -177 14530
rect -253 12730 -177 14270
rect -253 12470 -241 12730
rect -189 12470 -177 12730
rect -253 10930 -177 12470
rect -253 10670 -241 10930
rect -189 10670 -177 10930
rect -253 9130 -177 10670
rect -253 8870 -241 9130
rect -189 8870 -177 9130
rect -253 7330 -177 8870
rect -253 7070 -241 7330
rect -189 7070 -177 7330
rect -253 5530 -177 7070
rect -253 5270 -241 5530
rect -189 5270 -177 5530
rect -253 3730 -177 5270
rect -253 3470 -241 3730
rect -189 3470 -177 3730
rect -253 1930 -177 3470
rect -253 1670 -241 1930
rect -189 1670 -177 1930
rect -253 34 -177 1670
rect 23550 55933 23675 56012
rect 23550 55881 23587 55933
rect 23639 55881 23675 55933
rect 23550 55715 23675 55881
rect 23550 55663 23587 55715
rect 23639 55663 23675 55715
rect 23550 54133 23675 55663
rect 23550 54081 23587 54133
rect 23639 54081 23675 54133
rect 23550 53915 23675 54081
rect 23550 53863 23587 53915
rect 23639 53863 23675 53915
rect 23550 52333 23675 53863
rect 23550 52281 23587 52333
rect 23639 52281 23675 52333
rect 23550 52115 23675 52281
rect 23550 52063 23587 52115
rect 23639 52063 23675 52115
rect 23550 50533 23675 52063
rect 23550 50481 23587 50533
rect 23639 50481 23675 50533
rect 23550 50315 23675 50481
rect 23550 50263 23587 50315
rect 23639 50263 23675 50315
rect 23550 48733 23675 50263
rect 23550 48681 23587 48733
rect 23639 48681 23675 48733
rect 23550 48515 23675 48681
rect 23550 48463 23587 48515
rect 23639 48463 23675 48515
rect 23550 46933 23675 48463
rect 23550 46881 23587 46933
rect 23639 46881 23675 46933
rect 23550 46715 23675 46881
rect 23550 46663 23587 46715
rect 23639 46663 23675 46715
rect 23550 45133 23675 46663
rect 23550 45081 23587 45133
rect 23639 45081 23675 45133
rect 23550 44915 23675 45081
rect 23550 44863 23587 44915
rect 23639 44863 23675 44915
rect 23550 43333 23675 44863
rect 23550 43281 23587 43333
rect 23639 43281 23675 43333
rect 23550 43115 23675 43281
rect 23550 43063 23587 43115
rect 23639 43063 23675 43115
rect 23550 41533 23675 43063
rect 23550 41481 23587 41533
rect 23639 41481 23675 41533
rect 23550 41315 23675 41481
rect 23550 41263 23587 41315
rect 23639 41263 23675 41315
rect 23550 39733 23675 41263
rect 23550 39681 23587 39733
rect 23639 39681 23675 39733
rect 23550 39515 23675 39681
rect 23550 39463 23587 39515
rect 23639 39463 23675 39515
rect 23550 37933 23675 39463
rect 23550 37881 23587 37933
rect 23639 37881 23675 37933
rect 23550 37715 23675 37881
rect 23550 37663 23587 37715
rect 23639 37663 23675 37715
rect 23550 36133 23675 37663
rect 23550 36081 23587 36133
rect 23639 36081 23675 36133
rect 23550 35915 23675 36081
rect 23550 35863 23587 35915
rect 23639 35863 23675 35915
rect 23550 34333 23675 35863
rect 23550 34281 23587 34333
rect 23639 34281 23675 34333
rect 23550 34115 23675 34281
rect 23550 34063 23587 34115
rect 23639 34063 23675 34115
rect 23550 32533 23675 34063
rect 23550 32481 23587 32533
rect 23639 32481 23675 32533
rect 23550 32315 23675 32481
rect 23550 32263 23587 32315
rect 23639 32263 23675 32315
rect 23550 30733 23675 32263
rect 23550 30681 23587 30733
rect 23639 30681 23675 30733
rect 23550 30515 23675 30681
rect 23550 30463 23587 30515
rect 23639 30463 23675 30515
rect 23550 28933 23675 30463
rect 23550 28881 23587 28933
rect 23639 28881 23675 28933
rect 23550 28715 23675 28881
rect 23550 28663 23587 28715
rect 23639 28663 23675 28715
rect 23550 27133 23675 28663
rect 23550 27081 23587 27133
rect 23639 27081 23675 27133
rect 23550 26915 23675 27081
rect 23550 26863 23587 26915
rect 23639 26863 23675 26915
rect 23550 25337 23675 26863
rect 23550 25285 23587 25337
rect 23639 25285 23675 25337
rect 23550 25119 23675 25285
rect 23550 25067 23587 25119
rect 23639 25067 23675 25119
rect 23550 23533 23675 25067
rect 23550 23481 23587 23533
rect 23639 23481 23675 23533
rect 23550 23315 23675 23481
rect 23550 23263 23587 23315
rect 23639 23263 23675 23315
rect 23550 21737 23675 23263
rect 23550 21685 23587 21737
rect 23639 21685 23675 21737
rect 23550 21519 23675 21685
rect 23550 21467 23587 21519
rect 23639 21467 23675 21519
rect 23550 19933 23675 21467
rect 23550 19881 23587 19933
rect 23639 19881 23675 19933
rect 23550 19715 23675 19881
rect 23550 19663 23587 19715
rect 23639 19663 23675 19715
rect 23550 18137 23675 19663
rect 23550 18085 23587 18137
rect 23639 18085 23675 18137
rect 23550 17919 23675 18085
rect 23550 17867 23587 17919
rect 23639 17867 23675 17919
rect 23550 16333 23675 17867
rect 23550 16281 23587 16333
rect 23639 16281 23675 16333
rect 23550 16115 23675 16281
rect 23550 16063 23587 16115
rect 23639 16063 23675 16115
rect 23550 14537 23675 16063
rect 23550 14485 23587 14537
rect 23639 14485 23675 14537
rect 23550 14319 23675 14485
rect 23550 14267 23587 14319
rect 23639 14267 23675 14319
rect 23550 12733 23675 14267
rect 23550 12681 23587 12733
rect 23639 12681 23675 12733
rect 23550 12515 23675 12681
rect 23550 12463 23587 12515
rect 23639 12463 23675 12515
rect 23550 10937 23675 12463
rect 23550 10885 23587 10937
rect 23639 10885 23675 10937
rect 23550 10719 23675 10885
rect 23550 10667 23587 10719
rect 23639 10667 23675 10719
rect 23550 9133 23675 10667
rect 23550 9081 23587 9133
rect 23639 9081 23675 9133
rect 23550 8915 23675 9081
rect 23550 8863 23587 8915
rect 23639 8863 23675 8915
rect 23550 7337 23675 8863
rect 23550 7285 23587 7337
rect 23639 7285 23675 7337
rect 23550 7119 23675 7285
rect 23550 7067 23587 7119
rect 23639 7067 23675 7119
rect 23550 5533 23675 7067
rect 23550 5481 23587 5533
rect 23639 5481 23675 5533
rect 23550 5315 23675 5481
rect 23550 5263 23587 5315
rect 23639 5263 23675 5315
rect 23550 3737 23675 5263
rect 23550 3685 23587 3737
rect 23639 3685 23675 3737
rect 23550 3519 23675 3685
rect 23550 3467 23587 3519
rect 23639 3467 23675 3519
rect 23550 1933 23675 3467
rect 23550 1881 23587 1933
rect 23639 1881 23675 1933
rect 23550 1715 23675 1881
rect 23550 1663 23587 1715
rect 23639 1663 23675 1715
rect 23550 400 23675 1663
rect 23550 348 23587 400
rect 23639 348 23675 400
rect -358 24 -74 34
rect -358 -32 -348 24
rect -84 -32 -74 24
rect -358 -42 -74 -32
rect 22890 -857 23010 326
rect 22847 -955 23010 -857
rect 23190 -857 23310 326
rect 23550 182 23675 348
rect 23550 130 23587 182
rect 23639 130 23675 182
rect 23550 90 23675 130
rect 23190 -955 23318 -857
rect 22847 -1250 22903 -955
rect 23262 -1250 23318 -955
rect 23049 -25410 23179 -17598
<< via2 >>
rect -348 -32 -84 24
<< metal3 >>
rect -358 24 -74 72
rect -358 -32 -348 24
rect -84 -32 -74 24
rect -358 -68 -74 -32
rect 22329 -2910 23899 -1101
rect 22384 -8791 23899 -6814
rect 22279 -9117 23899 -8902
rect 22279 -9439 23899 -9223
rect 22279 -9760 23899 -9545
rect 22279 -10082 23899 -9867
rect 22279 -10774 23582 -10559
rect 22279 -11096 23582 -10881
rect 22279 -11418 23582 -11203
rect 22279 -11740 23582 -11524
rect 22384 -12288 23582 -11846
rect 22384 -13399 23899 -12944
rect 22426 -17210 23403 -14487
rect 22426 -20898 23403 -17496
rect 22351 -21764 23403 -21047
rect 22351 -23190 23403 -22379
rect 22426 -25051 23051 -23735
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_0
timestamp 1666464484
transform -1 0 600 0 1 11700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_1
timestamp 1666464484
transform -1 0 600 0 1 4500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_2
timestamp 1666464484
transform -1 0 600 0 1 8100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_3
timestamp 1666464484
transform -1 0 600 0 1 15300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_4
timestamp 1666464484
transform -1 0 600 0 1 9900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_5
timestamp 1666464484
transform -1 0 600 0 1 13500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_6
timestamp 1666464484
transform -1 0 600 0 1 2700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_7
timestamp 1666464484
transform -1 0 600 0 1 6300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_8
timestamp 1666464484
transform -1 0 600 0 1 900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_9
timestamp 1666464484
transform -1 0 600 0 1 29700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_10
timestamp 1666464484
transform -1 0 600 0 1 35100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_11
timestamp 1666464484
transform -1 0 600 0 1 33300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_12
timestamp 1666464484
transform -1 0 600 0 1 36900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_13
timestamp 1666464484
transform -1 0 600 0 1 31500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_14
timestamp 1666464484
transform -1 0 600 0 1 18900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_15
timestamp 1666464484
transform -1 0 600 0 1 26100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_16
timestamp 1666464484
transform -1 0 600 0 1 22500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_17
timestamp 1666464484
transform -1 0 600 0 1 24300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_18
timestamp 1666464484
transform -1 0 600 0 1 27900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_19
timestamp 1666464484
transform -1 0 600 0 1 20700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_20
timestamp 1666464484
transform -1 0 600 0 1 42300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_21
timestamp 1666464484
transform -1 0 600 0 1 45900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_22
timestamp 1666464484
transform -1 0 600 0 1 49500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_23
timestamp 1666464484
transform -1 0 600 0 1 56700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_24
timestamp 1666464484
transform -1 0 600 0 1 53100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_25
timestamp 1666464484
transform -1 0 600 0 1 40500
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_26
timestamp 1666464484
transform -1 0 600 0 1 44100
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_27
timestamp 1666464484
transform -1 0 600 0 1 47700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_28
timestamp 1666464484
transform -1 0 600 0 1 54900
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_29
timestamp 1666464484
transform -1 0 600 0 1 51300
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_30
timestamp 1666464484
transform -1 0 600 0 1 38700
box -68 -68 668 1868
use 018SRAM_cell1_2x_512x8m81  018SRAM_cell1_2x_512x8m81_31
timestamp 1666464484
transform -1 0 600 0 1 17100
box -68 -68 668 1868
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_0
timestamp 1666464484
transform -1 0 600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_512x8m81  018SRAM_cell1_512x8m81_1
timestamp 1666464484
transform -1 0 600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_0
timestamp 1666464484
transform -1 0 16800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_1
timestamp 1666464484
transform -1 0 16200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_2
timestamp 1666464484
transform -1 0 15600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_3
timestamp 1666464484
transform -1 0 15000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_4
timestamp 1666464484
transform -1 0 13800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_5
timestamp 1666464484
transform -1 0 14400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_6
timestamp 1666464484
transform -1 0 13200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_7
timestamp 1666464484
transform -1 0 12600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_8
timestamp 1666464484
transform -1 0 18000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_9
timestamp 1666464484
transform -1 0 18600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_10
timestamp 1666464484
transform -1 0 19800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_11
timestamp 1666464484
transform -1 0 19200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_12
timestamp 1666464484
transform -1 0 20400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_13
timestamp 1666464484
transform -1 0 21000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_14
timestamp 1666464484
transform -1 0 21600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_15
timestamp 1666464484
transform -1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_16
timestamp 1666464484
transform -1 0 7800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_17
timestamp 1666464484
transform -1 0 9000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_18
timestamp 1666464484
transform -1 0 8400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_19
timestamp 1666464484
transform -1 0 9600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_20
timestamp 1666464484
transform -1 0 10200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_21
timestamp 1666464484
transform -1 0 10800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_22
timestamp 1666464484
transform -1 0 11400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_23
timestamp 1666464484
transform -1 0 6000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_24
timestamp 1666464484
transform -1 0 5400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_25
timestamp 1666464484
transform -1 0 4800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_26
timestamp 1666464484
transform -1 0 4200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_27
timestamp 1666464484
transform -1 0 3000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_28
timestamp 1666464484
transform -1 0 3600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_29
timestamp 1666464484
transform -1 0 2400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_30
timestamp 1666464484
transform -1 0 1800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_31
timestamp 1666464484
transform -1 0 7200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_32
timestamp 1666464484
transform -1 0 4200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_33
timestamp 1666464484
transform -1 0 3000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_34
timestamp 1666464484
transform -1 0 3600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_35
timestamp 1666464484
transform -1 0 2400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_36
timestamp 1666464484
transform -1 0 1800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_37
timestamp 1666464484
transform -1 0 5400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_38
timestamp 1666464484
transform -1 0 4800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_39
timestamp 1666464484
transform -1 0 10800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_40
timestamp 1666464484
transform -1 0 7200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_41
timestamp 1666464484
transform -1 0 11400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_42
timestamp 1666464484
transform -1 0 7800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_43
timestamp 1666464484
transform -1 0 9000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_44
timestamp 1666464484
transform -1 0 8400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_45
timestamp 1666464484
transform -1 0 9600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_46
timestamp 1666464484
transform -1 0 10200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_47
timestamp 1666464484
transform -1 0 6000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_48
timestamp 1666464484
transform -1 0 13800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_49
timestamp 1666464484
transform -1 0 16200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_50
timestamp 1666464484
transform -1 0 12600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_51
timestamp 1666464484
transform -1 0 13200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_52
timestamp 1666464484
transform -1 0 16800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_53
timestamp 1666464484
transform -1 0 14400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_54
timestamp 1666464484
transform -1 0 15000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_55
timestamp 1666464484
transform -1 0 15600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_56
timestamp 1666464484
transform -1 0 19200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_57
timestamp 1666464484
transform -1 0 18600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_58
timestamp 1666464484
transform -1 0 21000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_59
timestamp 1666464484
transform -1 0 20400 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_60
timestamp 1666464484
transform -1 0 21600 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_61
timestamp 1666464484
transform -1 0 19800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_62
timestamp 1666464484
transform -1 0 22200 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_512x8m81  018SRAM_cell1_dummy_512x8m81_63
timestamp 1666464484
transform -1 0 18000 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_0
timestamp 1666464484
transform 1 0 22800 0 -1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_1
timestamp 1666464484
transform 1 0 22800 0 -1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_2
timestamp 1666464484
transform 1 0 22800 0 -1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_3
timestamp 1666464484
transform 1 0 22800 0 -1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_4
timestamp 1666464484
transform 1 0 22800 0 -1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_5
timestamp 1666464484
transform 1 0 22800 0 -1 18000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_6
timestamp 1666464484
transform 1 0 22800 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_7
timestamp 1666464484
transform 1 0 22800 0 -1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_8
timestamp 1666464484
transform 1 0 22800 0 -1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_9
timestamp 1666464484
transform 1 0 22800 0 -1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_10
timestamp 1666464484
transform 1 0 22800 0 1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_11
timestamp 1666464484
transform 1 0 22800 0 1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_12
timestamp 1666464484
transform 1 0 22800 0 1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_13
timestamp 1666464484
transform 1 0 22800 0 1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_14
timestamp 1666464484
transform 1 0 22800 0 1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_15
timestamp 1666464484
transform 1 0 22800 0 1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_16
timestamp 1666464484
transform 1 0 22800 0 1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_17
timestamp 1666464484
transform 1 0 22800 0 1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_18
timestamp 1666464484
transform 1 0 22800 0 1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_19
timestamp 1666464484
transform 1 0 22800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_20
timestamp 1666464484
transform 1 0 22800 0 -1 37800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_21
timestamp 1666464484
transform 1 0 22800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_22
timestamp 1666464484
transform 1 0 22800 0 -1 36000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_23
timestamp 1666464484
transform 1 0 22800 0 -1 34200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_24
timestamp 1666464484
transform 1 0 22800 0 -1 32400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_25
timestamp 1666464484
transform 1 0 22800 0 -1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_26
timestamp 1666464484
transform 1 0 22800 0 -1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_27
timestamp 1666464484
transform 1 0 22800 0 -1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_28
timestamp 1666464484
transform 1 0 22800 0 -1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_29
timestamp 1666464484
transform 1 0 22800 0 -1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_30
timestamp 1666464484
transform 1 0 22800 0 -1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_31
timestamp 1666464484
transform 1 0 22800 0 1 36000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_32
timestamp 1666464484
transform 1 0 22800 0 1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_33
timestamp 1666464484
transform 1 0 22800 0 1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_34
timestamp 1666464484
transform 1 0 22800 0 1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_35
timestamp 1666464484
transform 1 0 22800 0 1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_36
timestamp 1666464484
transform 1 0 22800 0 1 32400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_37
timestamp 1666464484
transform 1 0 22800 0 1 34200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_38
timestamp 1666464484
transform 1 0 22800 0 1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_39
timestamp 1666464484
transform 1 0 22800 0 1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_40
timestamp 1666464484
transform 1 0 22800 0 1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_41
timestamp 1666464484
transform 1 0 22800 0 1 37800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_42
timestamp 1666464484
transform 1 0 22800 0 -1 55800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_43
timestamp 1666464484
transform 1 0 22800 0 -1 52200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_44
timestamp 1666464484
transform 1 0 22800 0 -1 48600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_45
timestamp 1666464484
transform 1 0 22800 0 -1 43200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_46
timestamp 1666464484
transform 1 0 22800 0 -1 41400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_47
timestamp 1666464484
transform 1 0 22800 0 -1 57600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_48
timestamp 1666464484
transform 1 0 22800 0 -1 54000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_49
timestamp 1666464484
transform 1 0 22800 0 -1 50400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_50
timestamp 1666464484
transform 1 0 22800 0 -1 46800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_51
timestamp 1666464484
transform 1 0 22800 0 -1 45000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_52
timestamp 1666464484
transform 1 0 22800 0 -1 59400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_53
timestamp 1666464484
transform 1 0 22800 0 1 54000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_54
timestamp 1666464484
transform 1 0 22800 0 1 39600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_55
timestamp 1666464484
transform 1 0 22800 0 1 46800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_56
timestamp 1666464484
transform 1 0 22800 0 1 55800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_57
timestamp 1666464484
transform 1 0 22800 0 1 50400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_58
timestamp 1666464484
transform 1 0 22800 0 1 43200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_59
timestamp 1666464484
transform 1 0 22800 0 1 57600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_60
timestamp 1666464484
transform 1 0 22800 0 1 45000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_61
timestamp 1666464484
transform 1 0 22800 0 1 52200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_62
timestamp 1666464484
transform 1 0 22800 0 1 41400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_63
timestamp 1666464484
transform 1 0 22800 0 1 48600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_64
timestamp 1666464484
transform 1 0 22800 0 -1 39600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_512x8m81  018SRAM_cell1_dummy_R_512x8m81_65
timestamp 1666464484
transform 1 0 22800 0 1 18000
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_0
timestamp 1666464484
transform -1 0 17400 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_1
timestamp 1666464484
transform -1 0 6600 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_2
timestamp 1666464484
transform -1 0 1200 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_3
timestamp 1666464484
transform -1 0 6600 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_4
timestamp 1666464484
transform -1 0 17400 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_5
timestamp 1666464484
transform 1 0 22200 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_6
timestamp 1666464484
transform -1 0 12000 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_512x8m81  018SRAM_strap1_512x8m81_7
timestamp 1666464484
transform -1 0 12000 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_0
timestamp 1666464484
transform 1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_1
timestamp 1666464484
transform -1 0 1200 0 -1 3600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_2
timestamp 1666464484
transform -1 0 1200 0 -1 5400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_3
timestamp 1666464484
transform -1 0 1200 0 1 1800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_4
timestamp 1666464484
transform -1 0 1200 0 1 3600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_5
timestamp 1666464484
transform -1 0 1200 0 -1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_6
timestamp 1666464484
transform -1 0 1200 0 1 5400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_7
timestamp 1666464484
transform -1 0 1200 0 1 9000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_8
timestamp 1666464484
transform -1 0 1200 0 1 7200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_9
timestamp 1666464484
transform -1 0 1200 0 1 10800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_10
timestamp 1666464484
transform -1 0 1200 0 1 12600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_11
timestamp 1666464484
transform -1 0 1200 0 -1 1800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_12
timestamp 1666464484
transform -1 0 1200 0 -1 14400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_13
timestamp 1666464484
transform -1 0 1200 0 -1 18000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_14
timestamp 1666464484
transform -1 0 1200 0 -1 7200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_15
timestamp 1666464484
transform -1 0 1200 0 -1 10800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_16
timestamp 1666464484
transform -1 0 1200 0 1 14400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_17
timestamp 1666464484
transform -1 0 1200 0 -1 12600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_18
timestamp 1666464484
transform -1 0 1200 0 -1 9000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_19
timestamp 1666464484
transform -1 0 1200 0 1 16200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_20
timestamp 1666464484
transform -1 0 1200 0 1 34200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_21
timestamp 1666464484
transform -1 0 1200 0 1 36000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_22
timestamp 1666464484
transform -1 0 1200 0 1 37800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_23
timestamp 1666464484
transform -1 0 1200 0 -1 23400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_24
timestamp 1666464484
transform -1 0 1200 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_25
timestamp 1666464484
transform -1 0 1200 0 -1 36000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_26
timestamp 1666464484
transform -1 0 1200 0 -1 27000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_27
timestamp 1666464484
transform -1 0 1200 0 1 30600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_28
timestamp 1666464484
transform -1 0 1200 0 -1 28800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_29
timestamp 1666464484
transform -1 0 1200 0 -1 34200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_30
timestamp 1666464484
transform -1 0 1200 0 -1 32400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_31
timestamp 1666464484
transform -1 0 1200 0 1 27000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_32
timestamp 1666464484
transform -1 0 1200 0 -1 37800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_33
timestamp 1666464484
transform -1 0 1200 0 1 28800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_34
timestamp 1666464484
transform -1 0 1200 0 -1 19800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_35
timestamp 1666464484
transform -1 0 1200 0 1 23400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_36
timestamp 1666464484
transform -1 0 1200 0 1 25200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_37
timestamp 1666464484
transform -1 0 1200 0 1 21600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_38
timestamp 1666464484
transform -1 0 1200 0 1 19800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_39
timestamp 1666464484
transform -1 0 1200 0 -1 25200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_40
timestamp 1666464484
transform -1 0 1200 0 1 32400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_41
timestamp 1666464484
transform -1 0 1200 0 -1 21600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_42
timestamp 1666464484
transform -1 0 1200 0 -1 50400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_43
timestamp 1666464484
transform -1 0 1200 0 1 57600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_44
timestamp 1666464484
transform -1 0 1200 0 1 54000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_45
timestamp 1666464484
transform -1 0 1200 0 1 46800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_46
timestamp 1666464484
transform -1 0 1200 0 1 41400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_47
timestamp 1666464484
transform -1 0 1200 0 1 39600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_48
timestamp 1666464484
transform -1 0 1200 0 1 43200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_49
timestamp 1666464484
transform -1 0 1200 0 1 45000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_50
timestamp 1666464484
transform -1 0 1200 0 1 55800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_51
timestamp 1666464484
transform -1 0 1200 0 1 52200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_52
timestamp 1666464484
transform -1 0 1200 0 1 50400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_53
timestamp 1666464484
transform -1 0 1200 0 1 48600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_54
timestamp 1666464484
transform -1 0 1200 0 -1 59400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_55
timestamp 1666464484
transform -1 0 1200 0 -1 46800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_56
timestamp 1666464484
transform -1 0 1200 0 -1 57600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_57
timestamp 1666464484
transform -1 0 1200 0 -1 45000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_58
timestamp 1666464484
transform -1 0 1200 0 -1 52200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_59
timestamp 1666464484
transform -1 0 1200 0 -1 48600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_60
timestamp 1666464484
transform -1 0 1200 0 -1 54000
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_61
timestamp 1666464484
transform -1 0 1200 0 -1 41400
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_62
timestamp 1666464484
transform -1 0 1200 0 -1 43200
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_63
timestamp 1666464484
transform -1 0 1200 0 -1 55800
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_64
timestamp 1666464484
transform -1 0 1200 0 -1 39600
box -68 -68 668 968
use 018SRAM_strap1_bndry_512x8m81  018SRAM_strap1_bndry_512x8m81_65
timestamp 1666464484
transform -1 0 1200 0 1 18000
box -68 -68 668 968
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_0
timestamp 1666464484
transform 1 0 23318 0 1 -22942
box 0 0 1 1
use M1_NWELL$$44998700_512x8m81  M1_NWELL$$44998700_512x8m81_1
timestamp 1666464484
transform 1 0 22774 0 1 -22942
box 0 0 1 1
use M1_NWELL$$46277676_512x8m81  M1_NWELL$$46277676_512x8m81_0
timestamp 1666464484
transform 1 0 23050 0 1 -14622
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_0
timestamp 1666464484
transform 1 0 23615 0 -1 7200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_1
timestamp 1666464484
transform 1 0 23615 0 -1 5400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_2
timestamp 1666464484
transform 1 0 23615 0 -1 1800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_3
timestamp 1666464484
transform 1 0 23615 0 -1 240
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_4
timestamp 1666464484
transform 1 0 23615 0 -1 16200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_5
timestamp 1666464484
transform 1 0 23615 0 -1 12600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_6
timestamp 1666464484
transform 1 0 23615 0 -1 9000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_7
timestamp 1666464484
transform 1 0 23615 0 -1 14400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_8
timestamp 1666464484
transform 1 0 23615 0 -1 10800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_9
timestamp 1666464484
transform 1 0 23615 0 -1 3600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_10
timestamp 1666464484
transform 1 0 23615 0 -1 21600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_11
timestamp 1666464484
transform 1 0 23615 0 -1 37800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_12
timestamp 1666464484
transform 1 0 23615 0 -1 36000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_13
timestamp 1666464484
transform 1 0 23615 0 -1 34200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_14
timestamp 1666464484
transform 1 0 23615 0 -1 32400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_15
timestamp 1666464484
transform 1 0 23615 0 -1 30600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_16
timestamp 1666464484
transform 1 0 23615 0 -1 27000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_17
timestamp 1666464484
transform 1 0 23615 0 -1 23400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_18
timestamp 1666464484
transform 1 0 23615 0 -1 19800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_19
timestamp 1666464484
transform 1 0 23615 0 -1 28800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_20
timestamp 1666464484
transform 1 0 23615 0 -1 25200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_21
timestamp 1666464484
transform 1 0 23615 0 -1 55800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_22
timestamp 1666464484
transform 1 0 23615 0 -1 54000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_23
timestamp 1666464484
transform 1 0 23615 0 -1 52200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_24
timestamp 1666464484
transform 1 0 23615 0 -1 50400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_25
timestamp 1666464484
transform 1 0 23615 0 -1 48600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_26
timestamp 1666464484
transform 1 0 23615 0 -1 46800
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_27
timestamp 1666464484
transform 1 0 23615 0 -1 45000
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_28
timestamp 1666464484
transform 1 0 23615 0 -1 43200
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_29
timestamp 1666464484
transform 1 0 23615 0 -1 41400
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_30
timestamp 1666464484
transform 1 0 23615 0 -1 39600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_31
timestamp 1666464484
transform 1 0 23615 0 -1 57600
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_32
timestamp 1666464484
transform 1 0 23615 0 -1 59160
box 0 0 1 1
use M1_POLY2$$44754988_512x8m81  M1_POLY2$$44754988_512x8m81_33
timestamp 1666464484
transform 1 0 23615 0 -1 18000
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_0
timestamp 1666464484
transform -1 0 22809 0 1 -19544
box 0 0 1 1
use M1_POLY2$$46559276_512x8m81_0  M1_POLY2$$46559276_512x8m81_0_1
timestamp 1666464484
transform 1 0 23393 0 1 -15883
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_0
timestamp 1666464484
transform 1 0 -215 0 1 141
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_1
timestamp 1666464484
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_2
timestamp 1666464484
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_3
timestamp 1666464484
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_4
timestamp 1666464484
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_5
timestamp 1666464484
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_6
timestamp 1666464484
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_7
timestamp 1666464484
transform 1 0 -215 0 1 16200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_8
timestamp 1666464484
transform 1 0 -215 0 1 18000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_9
timestamp 1666464484
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_10
timestamp 1666464484
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_11
timestamp 1666464484
transform 1 0 -215 0 1 21600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_12
timestamp 1666464484
transform 1 0 -215 0 1 19800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_13
timestamp 1666464484
transform 1 0 -215 0 1 23400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_14
timestamp 1666464484
transform 1 0 -215 0 1 25200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_15
timestamp 1666464484
transform 1 0 -215 0 1 28800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_16
timestamp 1666464484
transform 1 0 -215 0 1 27000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_17
timestamp 1666464484
transform 1 0 -215 0 1 30600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_18
timestamp 1666464484
transform 1 0 -215 0 1 32400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_19
timestamp 1666464484
transform 1 0 -215 0 1 36000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_20
timestamp 1666464484
transform 1 0 -215 0 1 34200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_21
timestamp 1666464484
transform 1 0 -215 0 1 37800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_22
timestamp 1666464484
transform 1 0 -215 0 1 39600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_23
timestamp 1666464484
transform 1 0 -215 0 1 43200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_24
timestamp 1666464484
transform 1 0 -215 0 1 41400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_25
timestamp 1666464484
transform 1 0 -215 0 1 45000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_26
timestamp 1666464484
transform 1 0 -215 0 1 46800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_27
timestamp 1666464484
transform 1 0 -215 0 1 50400
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_28
timestamp 1666464484
transform 1 0 -215 0 1 48600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_29
timestamp 1666464484
transform 1 0 -215 0 1 52200
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_30
timestamp 1666464484
transform 1 0 -215 0 1 54000
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_31
timestamp 1666464484
transform 1 0 -215 0 1 57600
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_32
timestamp 1666464484
transform 1 0 -215 0 1 55800
box 0 0 1 1
use M1_POLY24310591302019_512x8m81  M1_POLY24310591302019_512x8m81_33
timestamp 1666464484
transform 1 0 -215 0 1 59259
box 0 0 1 1
use M1_PSUB$$46274604_512x8m81  M1_PSUB$$46274604_512x8m81_0
timestamp 1666464484
transform 1 0 23107 0 1 -16617
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_0
timestamp 1666464484
transform 1 0 23613 0 -1 16198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_1
timestamp 1666464484
transform 1 0 23613 0 -1 12598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_2
timestamp 1666464484
transform 1 0 23613 0 -1 8998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_3
timestamp 1666464484
transform 1 0 23613 0 -1 5398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_4
timestamp 1666464484
transform 1 0 23613 0 -1 1798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_5
timestamp 1666464484
transform 1 0 23613 0 -1 10802
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_6
timestamp 1666464484
transform 1 0 23613 0 -1 3602
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_7
timestamp 1666464484
transform 1 0 23613 0 -1 265
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_8
timestamp 1666464484
transform 1 0 23613 0 -1 14402
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_9
timestamp 1666464484
transform 1 0 23613 0 -1 7202
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_10
timestamp 1666464484
transform 1 0 23613 0 -1 32398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_11
timestamp 1666464484
transform 1 0 23613 0 -1 30598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_12
timestamp 1666464484
transform 1 0 23613 0 -1 26998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_13
timestamp 1666464484
transform 1 0 23613 0 -1 23398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_14
timestamp 1666464484
transform 1 0 23613 0 -1 19798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_15
timestamp 1666464484
transform 1 0 23613 0 -1 25202
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_16
timestamp 1666464484
transform 1 0 23613 0 -1 28798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_17
timestamp 1666464484
transform 1 0 23613 0 -1 37798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_18
timestamp 1666464484
transform 1 0 23613 0 -1 21602
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_19
timestamp 1666464484
transform 1 0 23613 0 -1 35998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_20
timestamp 1666464484
transform 1 0 23613 0 -1 34198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_21
timestamp 1666464484
transform 1 0 23613 0 -1 55798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_22
timestamp 1666464484
transform 1 0 23613 0 -1 53998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_23
timestamp 1666464484
transform 1 0 23613 0 -1 52198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_24
timestamp 1666464484
transform 1 0 23613 0 -1 50398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_25
timestamp 1666464484
transform 1 0 23613 0 -1 48598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_26
timestamp 1666464484
transform 1 0 23613 0 -1 46798
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_27
timestamp 1666464484
transform 1 0 23613 0 -1 44998
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_28
timestamp 1666464484
transform 1 0 23613 0 -1 43198
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_29
timestamp 1666464484
transform 1 0 23613 0 -1 41398
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_30
timestamp 1666464484
transform 1 0 23613 0 -1 39598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_31
timestamp 1666464484
transform 1 0 23613 0 -1 59135
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_32
timestamp 1666464484
transform 1 0 23613 0 -1 57598
box 0 0 1 1
use M2_M1$$43375660_512x8m81  M2_M1$$43375660_512x8m81_33
timestamp 1666464484
transform 1 0 23613 0 -1 18002
box 0 0 1 1
use M2_M1$$47117356_512x8m81  M2_M1$$47117356_512x8m81_0
timestamp 1666464484
transform 1 0 23114 0 1 -20269
box -65 -2678 65 2678
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_0
timestamp 1666464484
transform 1 0 -215 0 1 1800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_1
timestamp 1666464484
transform 1 0 -215 0 1 3600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_2
timestamp 1666464484
transform 1 0 -215 0 1 5400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_3
timestamp 1666464484
transform 1 0 -215 0 1 7200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_4
timestamp 1666464484
transform 1 0 -215 0 1 9000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_5
timestamp 1666464484
transform 1 0 -215 0 1 10800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_6
timestamp 1666464484
transform 1 0 -215 0 1 12600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_7
timestamp 1666464484
transform 1 0 -215 0 1 14400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_8
timestamp 1666464484
transform 1 0 -215 0 1 16200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_9
timestamp 1666464484
transform 1 0 -215 0 1 18000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_10
timestamp 1666464484
transform 1 0 -215 0 1 37800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_11
timestamp 1666464484
transform 1 0 -215 0 1 36000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_12
timestamp 1666464484
transform 1 0 -215 0 1 34200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_13
timestamp 1666464484
transform 1 0 -215 0 1 32400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_14
timestamp 1666464484
transform 1 0 -215 0 1 30600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_15
timestamp 1666464484
transform 1 0 -215 0 1 28800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_16
timestamp 1666464484
transform 1 0 -215 0 1 27000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_17
timestamp 1666464484
transform 1 0 -215 0 1 25200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_18
timestamp 1666464484
transform 1 0 -215 0 1 19800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_19
timestamp 1666464484
transform 1 0 -215 0 1 21600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_20
timestamp 1666464484
transform 1 0 -219 0 1 23400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_21
timestamp 1666464484
transform 1 0 -215 0 1 57599
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_22
timestamp 1666464484
transform 1 0 -215 0 1 55800
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_23
timestamp 1666464484
transform 1 0 -215 0 1 54000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_24
timestamp 1666464484
transform 1 0 -215 0 1 52200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_25
timestamp 1666464484
transform 1 0 -215 0 1 50399
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_26
timestamp 1666464484
transform 1 0 -215 0 1 48600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_27
timestamp 1666464484
transform 1 0 -215 0 1 46801
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_28
timestamp 1666464484
transform 1 0 -215 0 1 45000
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_29
timestamp 1666464484
transform 1 0 -215 0 1 43200
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_30
timestamp 1666464484
transform 1 0 -215 0 1 41400
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_31
timestamp 1666464484
transform 1 0 -215 0 1 39600
box 0 0 1 1
use M2_M14310591302018_512x8m81  M2_M14310591302018_512x8m81_32
timestamp 1666464484
transform 1 0 -215 0 1 59198
box 0 0 1 1
use M3_M24310591302029_512x8m81  M3_M24310591302029_512x8m81_0
timestamp 1666464484
transform 0 -1 -216 1 0 -4
box 0 0 1 1
use nmos_5p04310591302096_512x8m81  nmos_5p04310591302096_512x8m81_0
timestamp 1666464484
transform 1 0 22940 0 1 -19403
box -88 -44 432 1744
use nmos_5p04310591302098_512x8m81  nmos_5p04310591302098_512x8m81_0
timestamp 1666464484
transform 1 0 22936 0 1 -16318
box -88 -44 432 320
use pmos_5p04310591302095_512x8m81  pmos_5p04310591302095_512x8m81_0
timestamp 1666464484
transform 1 0 22936 0 1 -15738
box -208 -120 552 822
use pmos_5p04310591302097_512x8m81  pmos_5p04310591302097_512x8m81_0
timestamp 1666464484
transform 1 0 22940 0 -1 -19684
box -208 -120 552 2248
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_0
timestamp 1666464484
transform 1 0 23283 0 1 -18447
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_1
timestamp 1666464484
transform 1 0 23285 0 1 -15470
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_2
timestamp 1666464484
transform 1 0 23288 0 1 -22897
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_3
timestamp 1666464484
transform 1 0 22846 0 1 -22711
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_4
timestamp 1666464484
transform 1 0 22842 0 1 -17909
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_5
timestamp 1666464484
transform 1 0 22842 0 1 -19052
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_6
timestamp 1666464484
transform 1 0 22837 0 1 -15470
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_7
timestamp 1666464484
transform 1 0 23288 0 1 -22711
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_8
timestamp 1666464484
transform 1 0 22842 0 1 -18447
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_9
timestamp 1666464484
transform 1 0 22846 0 1 -22897
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_10
timestamp 1666464484
transform 1 0 23283 0 1 -17909
box 0 -1 93 308
use via1_2_x2_512x8m81_0  via1_2_x2_512x8m81_0_11
timestamp 1666464484
transform 1 0 23283 0 1 -19052
box 0 -1 93 308
use via1_2_x2_R90_512x8m81_0  via1_2_x2_R90_512x8m81_0_0
timestamp 1666464484
transform 0 -1 23187 1 0 -14670
box 0 -1 93 308
use via1_2_x2_R270_512x8m81_0  via1_2_x2_R270_512x8m81_0_0
timestamp 1666464484
transform 0 1 22794 -1 0 -12002
box -1 -1 96 308
use ypass_gate_512x8m81_0  ypass_gate_512x8m81_0_0
timestamp 1666464484
transform -1 0 23395 0 1 -13448
box -221 -1 930 12370
<< labels >>
rlabel metal2 s 902 880 902 880 4 VDD
rlabel metal3 s 22866 1818 22866 1818 4 VSS
rlabel metal3 s 534 1818 534 1818 4 VSS
rlabel metal3 s 22866 893 22866 893 4 VDD
rlabel metal3 s 534 893 534 893 4 VDD
rlabel metal3 s 534 29693 534 29693 4 VDD
rlabel metal3 s 162 58942 162 58942 4 DWL
rlabel metal3 s 534 30618 534 30618 4 VSS
rlabel metal3 s 22541 -21185 22541 -21185 4 vdd
port 1 nsew
rlabel metal3 s 22541 -14704 22541 -14704 4 vdd
port 1 nsew
rlabel metal3 s 22644 -13162 22644 -13162 4 vss
port 2 nsew
rlabel metal3 s 22541 -12038 22541 -12038 4 vdd
port 1 nsew
rlabel metal3 s 22541 -6717 22541 -6717 4 vss
port 2 nsew
rlabel metal3 s 22541 -1276 22541 -1276 4 vdd
port 1 nsew
rlabel metal1 s 23127 -25252 23127 -25252 4 tblhl
port 3 nsew
rlabel metal1 s 23039 -16606 23039 -16606 4 vss
port 2 nsew
rlabel metal1 s 23037 -3126 23037 -3126 4 pcb
port 4 nsew
rlabel metal1 s 23037 -3126 23037 -3126 4 pcb
port 4 nsew
<< properties >>
string GDS_END 2520116
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2481544
<< end >>
