magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 178
rect 224 0 344 178
rect 448 0 568 178
rect 672 0 792 178
rect 896 0 1016 178
rect 1120 0 1240 178
rect 1344 0 1464 178
<< mvndiff >>
rect -88 165 0 178
rect -88 119 -75 165
rect -29 119 0 165
rect -88 59 0 119
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 165 224 178
rect 120 119 149 165
rect 195 119 224 165
rect 120 59 224 119
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 165 448 178
rect 344 119 373 165
rect 419 119 448 165
rect 344 59 448 119
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 165 672 178
rect 568 119 597 165
rect 643 119 672 165
rect 568 59 672 119
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 165 896 178
rect 792 119 821 165
rect 867 119 896 165
rect 792 59 896 119
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 165 1120 178
rect 1016 119 1045 165
rect 1091 119 1120 165
rect 1016 59 1120 119
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 165 1344 178
rect 1240 119 1269 165
rect 1315 119 1344 165
rect 1240 59 1344 119
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 165 1552 178
rect 1464 119 1493 165
rect 1539 119 1552 165
rect 1464 59 1552 119
rect 1464 13 1493 59
rect 1539 13 1552 59
rect 1464 0 1552 13
<< mvndiffc >>
rect -75 119 -29 165
rect -75 13 -29 59
rect 149 119 195 165
rect 149 13 195 59
rect 373 119 419 165
rect 373 13 419 59
rect 597 119 643 165
rect 597 13 643 59
rect 821 119 867 165
rect 821 13 867 59
rect 1045 119 1091 165
rect 1045 13 1091 59
rect 1269 119 1315 165
rect 1269 13 1315 59
rect 1493 119 1539 165
rect 1493 13 1539 59
<< polysilicon >>
rect 0 178 120 222
rect 224 178 344 222
rect 448 178 568 222
rect 672 178 792 222
rect 896 178 1016 222
rect 1120 178 1240 222
rect 1344 178 1464 222
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
<< metal1 >>
rect -75 165 -29 178
rect -75 59 -29 119
rect -75 0 -29 13
rect 149 165 195 178
rect 149 59 195 119
rect 149 0 195 13
rect 373 165 419 178
rect 373 59 419 119
rect 373 0 419 13
rect 597 165 643 178
rect 597 59 643 119
rect 597 0 643 13
rect 821 165 867 178
rect 821 59 867 119
rect 821 0 867 13
rect 1045 165 1091 178
rect 1045 59 1091 119
rect 1045 0 1091 13
rect 1269 165 1315 178
rect 1269 59 1315 119
rect 1269 0 1315 13
rect 1493 165 1539 178
rect 1493 59 1539 119
rect 1493 0 1539 13
<< labels >>
flabel metal1 s -52 89 -52 89 0 FreeSans 200 0 0 0 S
flabel metal1 s 1516 89 1516 89 0 FreeSans 200 0 0 0 D
flabel metal1 s 172 89 172 89 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 89 396 89 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 89 620 89 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 89 844 89 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 89 1068 89 0 FreeSans 200 0 0 0 D
flabel metal1 s 1292 89 1292 89 0 FreeSans 200 0 0 0 S
<< properties >>
string GDS_END 568274
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 564062
<< end >>
