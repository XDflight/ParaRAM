magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 2268
<< mvndiff >>
rect -88 2255 0 2268
rect -88 2209 -75 2255
rect -29 2209 0 2255
rect -88 2151 0 2209
rect -88 2105 -75 2151
rect -29 2105 0 2151
rect -88 2047 0 2105
rect -88 2001 -75 2047
rect -29 2001 0 2047
rect -88 1943 0 2001
rect -88 1897 -75 1943
rect -29 1897 0 1943
rect -88 1839 0 1897
rect -88 1793 -75 1839
rect -29 1793 0 1839
rect -88 1735 0 1793
rect -88 1689 -75 1735
rect -29 1689 0 1735
rect -88 1631 0 1689
rect -88 1585 -75 1631
rect -29 1585 0 1631
rect -88 1527 0 1585
rect -88 1481 -75 1527
rect -29 1481 0 1527
rect -88 1423 0 1481
rect -88 1377 -75 1423
rect -29 1377 0 1423
rect -88 1319 0 1377
rect -88 1273 -75 1319
rect -29 1273 0 1319
rect -88 1214 0 1273
rect -88 1168 -75 1214
rect -29 1168 0 1214
rect -88 1109 0 1168
rect -88 1063 -75 1109
rect -29 1063 0 1109
rect -88 1004 0 1063
rect -88 958 -75 1004
rect -29 958 0 1004
rect -88 899 0 958
rect -88 853 -75 899
rect -29 853 0 899
rect -88 794 0 853
rect -88 748 -75 794
rect -29 748 0 794
rect -88 689 0 748
rect -88 643 -75 689
rect -29 643 0 689
rect -88 584 0 643
rect -88 538 -75 584
rect -29 538 0 584
rect -88 479 0 538
rect -88 433 -75 479
rect -29 433 0 479
rect -88 374 0 433
rect -88 328 -75 374
rect -29 328 0 374
rect -88 269 0 328
rect -88 223 -75 269
rect -29 223 0 269
rect -88 164 0 223
rect -88 118 -75 164
rect -29 118 0 164
rect -88 59 0 118
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 2255 208 2268
rect 120 2209 149 2255
rect 195 2209 208 2255
rect 120 2151 208 2209
rect 120 2105 149 2151
rect 195 2105 208 2151
rect 120 2047 208 2105
rect 120 2001 149 2047
rect 195 2001 208 2047
rect 120 1943 208 2001
rect 120 1897 149 1943
rect 195 1897 208 1943
rect 120 1839 208 1897
rect 120 1793 149 1839
rect 195 1793 208 1839
rect 120 1735 208 1793
rect 120 1689 149 1735
rect 195 1689 208 1735
rect 120 1631 208 1689
rect 120 1585 149 1631
rect 195 1585 208 1631
rect 120 1527 208 1585
rect 120 1481 149 1527
rect 195 1481 208 1527
rect 120 1423 208 1481
rect 120 1377 149 1423
rect 195 1377 208 1423
rect 120 1319 208 1377
rect 120 1273 149 1319
rect 195 1273 208 1319
rect 120 1214 208 1273
rect 120 1168 149 1214
rect 195 1168 208 1214
rect 120 1109 208 1168
rect 120 1063 149 1109
rect 195 1063 208 1109
rect 120 1004 208 1063
rect 120 958 149 1004
rect 195 958 208 1004
rect 120 899 208 958
rect 120 853 149 899
rect 195 853 208 899
rect 120 794 208 853
rect 120 748 149 794
rect 195 748 208 794
rect 120 689 208 748
rect 120 643 149 689
rect 195 643 208 689
rect 120 584 208 643
rect 120 538 149 584
rect 195 538 208 584
rect 120 479 208 538
rect 120 433 149 479
rect 195 433 208 479
rect 120 374 208 433
rect 120 328 149 374
rect 195 328 208 374
rect 120 269 208 328
rect 120 223 149 269
rect 195 223 208 269
rect 120 164 208 223
rect 120 118 149 164
rect 195 118 208 164
rect 120 59 208 118
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 2209 -29 2255
rect -75 2105 -29 2151
rect -75 2001 -29 2047
rect -75 1897 -29 1943
rect -75 1793 -29 1839
rect -75 1689 -29 1735
rect -75 1585 -29 1631
rect -75 1481 -29 1527
rect -75 1377 -29 1423
rect -75 1273 -29 1319
rect -75 1168 -29 1214
rect -75 1063 -29 1109
rect -75 958 -29 1004
rect -75 853 -29 899
rect -75 748 -29 794
rect -75 643 -29 689
rect -75 538 -29 584
rect -75 433 -29 479
rect -75 328 -29 374
rect -75 223 -29 269
rect -75 118 -29 164
rect -75 13 -29 59
rect 149 2209 195 2255
rect 149 2105 195 2151
rect 149 2001 195 2047
rect 149 1897 195 1943
rect 149 1793 195 1839
rect 149 1689 195 1735
rect 149 1585 195 1631
rect 149 1481 195 1527
rect 149 1377 195 1423
rect 149 1273 195 1319
rect 149 1168 195 1214
rect 149 1063 195 1109
rect 149 958 195 1004
rect 149 853 195 899
rect 149 748 195 794
rect 149 643 195 689
rect 149 538 195 584
rect 149 433 195 479
rect 149 328 195 374
rect 149 223 195 269
rect 149 118 195 164
rect 149 13 195 59
<< polysilicon >>
rect 0 2268 120 2312
rect 0 -44 120 0
<< metal1 >>
rect -75 2255 -29 2268
rect -75 2151 -29 2209
rect -75 2047 -29 2105
rect -75 1943 -29 2001
rect -75 1839 -29 1897
rect -75 1735 -29 1793
rect -75 1631 -29 1689
rect -75 1527 -29 1585
rect -75 1423 -29 1481
rect -75 1319 -29 1377
rect -75 1214 -29 1273
rect -75 1109 -29 1168
rect -75 1004 -29 1063
rect -75 899 -29 958
rect -75 794 -29 853
rect -75 689 -29 748
rect -75 584 -29 643
rect -75 479 -29 538
rect -75 374 -29 433
rect -75 269 -29 328
rect -75 164 -29 223
rect -75 59 -29 118
rect -75 0 -29 13
rect 149 2255 195 2268
rect 149 2151 195 2209
rect 149 2047 195 2105
rect 149 1943 195 2001
rect 149 1839 195 1897
rect 149 1735 195 1793
rect 149 1631 195 1689
rect 149 1527 195 1585
rect 149 1423 195 1481
rect 149 1319 195 1377
rect 149 1214 195 1273
rect 149 1109 195 1168
rect 149 1004 195 1063
rect 149 899 195 958
rect 149 794 195 853
rect 149 689 195 748
rect 149 584 195 643
rect 149 479 195 538
rect 149 374 195 433
rect 149 269 195 328
rect 149 164 195 223
rect 149 59 195 118
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1134 -52 1134 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 1134 172 1134 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 116212
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 112500
<< end >>
