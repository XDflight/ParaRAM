magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 3222 1094
<< pwell >>
rect -86 -86 3222 453
<< mvnmos >>
rect 124 156 244 296
rect 348 156 468 296
rect 572 156 692 296
rect 796 156 916 296
rect 975 156 1095 296
rect 1199 156 1319 296
rect 1655 137 1775 277
rect 1879 137 1999 277
rect 2247 122 2367 322
rect 2415 122 2535 322
rect 2639 122 2759 322
rect 2863 122 2983 322
<< mvpmos >>
rect 214 576 314 852
rect 362 576 462 852
rect 582 576 682 852
rect 884 576 984 852
rect 1032 576 1132 852
rect 1236 576 1336 852
rect 1615 573 1715 849
rect 1819 573 1919 849
rect 2257 573 2357 939
rect 2461 573 2561 939
rect 2665 573 2765 939
rect 2869 573 2969 939
<< mvndiff >>
rect 36 215 124 296
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 296
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 215 572 296
rect 468 169 497 215
rect 543 169 572 215
rect 468 156 572 169
rect 692 215 796 296
rect 692 169 721 215
rect 767 169 796 215
rect 692 156 796 169
rect 916 156 975 296
rect 1095 215 1199 296
rect 1095 169 1124 215
rect 1170 169 1199 215
rect 1095 156 1199 169
rect 1319 215 1407 296
rect 1319 169 1348 215
rect 1394 169 1407 215
rect 1319 156 1407 169
rect 2159 309 2247 322
rect 1567 215 1655 277
rect 1567 169 1580 215
rect 1626 169 1655 215
rect 1567 137 1655 169
rect 1775 215 1879 277
rect 1775 169 1804 215
rect 1850 169 1879 215
rect 1775 137 1879 169
rect 1999 196 2087 277
rect 1999 150 2028 196
rect 2074 150 2087 196
rect 1999 137 2087 150
rect 2159 169 2172 309
rect 2218 169 2247 309
rect 2159 122 2247 169
rect 2367 122 2415 322
rect 2535 275 2639 322
rect 2535 135 2564 275
rect 2610 135 2639 275
rect 2535 122 2639 135
rect 2759 309 2863 322
rect 2759 169 2788 309
rect 2834 169 2863 309
rect 2759 122 2863 169
rect 2983 275 3071 322
rect 2983 135 3012 275
rect 3058 135 3071 275
rect 2983 122 3071 135
<< mvpdiff >>
rect 126 839 214 852
rect 126 699 139 839
rect 185 699 214 839
rect 126 576 214 699
rect 314 576 362 852
rect 462 576 582 852
rect 682 839 884 852
rect 682 699 711 839
rect 757 699 884 839
rect 682 576 884 699
rect 984 576 1032 852
rect 1132 827 1236 852
rect 1132 781 1161 827
rect 1207 781 1236 827
rect 1132 576 1236 781
rect 1336 839 1424 852
rect 1336 699 1365 839
rect 1411 699 1424 839
rect 1336 576 1424 699
rect 1527 632 1615 849
rect 1527 586 1540 632
rect 1586 586 1615 632
rect 1527 573 1615 586
rect 1715 827 1819 849
rect 1715 781 1744 827
rect 1790 781 1819 827
rect 1715 573 1819 781
rect 1919 632 2007 849
rect 1919 586 1948 632
rect 1994 586 2007 632
rect 1919 573 2007 586
rect 2169 827 2257 939
rect 2169 781 2182 827
rect 2228 781 2257 827
rect 2169 573 2257 781
rect 2357 726 2461 939
rect 2357 586 2386 726
rect 2432 586 2461 726
rect 2357 573 2461 586
rect 2561 839 2665 939
rect 2561 699 2590 839
rect 2636 699 2665 839
rect 2561 573 2665 699
rect 2765 726 2869 939
rect 2765 586 2794 726
rect 2840 586 2869 726
rect 2765 573 2869 586
rect 2969 839 3057 939
rect 2969 699 2998 839
rect 3044 699 3057 839
rect 2969 573 3057 699
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 497 169 543 215
rect 721 169 767 215
rect 1124 169 1170 215
rect 1348 169 1394 215
rect 1580 169 1626 215
rect 1804 169 1850 215
rect 2028 150 2074 196
rect 2172 169 2218 309
rect 2564 135 2610 275
rect 2788 169 2834 309
rect 3012 135 3058 275
<< mvpdiffc >>
rect 139 699 185 839
rect 711 699 757 839
rect 1161 781 1207 827
rect 1365 699 1411 839
rect 1540 586 1586 632
rect 1744 781 1790 827
rect 1948 586 1994 632
rect 2182 781 2228 827
rect 2386 586 2432 726
rect 2590 699 2636 839
rect 2794 586 2840 726
rect 2998 699 3044 839
<< polysilicon >>
rect 884 944 1715 984
rect 214 852 314 896
rect 362 852 462 896
rect 582 852 682 896
rect 884 852 984 944
rect 1032 852 1132 896
rect 1236 852 1336 896
rect 1615 849 1715 944
rect 2257 939 2357 983
rect 2461 939 2561 983
rect 2665 939 2765 983
rect 2869 939 2969 983
rect 1819 849 1919 893
rect 214 532 314 576
rect 214 483 254 532
rect 362 483 462 576
rect 124 470 254 483
rect 124 424 142 470
rect 188 456 254 470
rect 348 470 462 483
rect 582 516 682 576
rect 884 543 984 576
rect 582 476 836 516
rect 884 497 897 543
rect 943 497 984 543
rect 884 484 984 497
rect 188 424 244 456
rect 124 296 244 424
rect 348 424 361 470
rect 407 424 462 470
rect 348 340 462 424
rect 572 415 748 428
rect 572 369 689 415
rect 735 369 748 415
rect 572 356 748 369
rect 348 296 468 340
rect 572 296 692 356
rect 796 340 836 476
rect 1032 483 1132 576
rect 1236 532 1336 576
rect 1236 483 1319 532
rect 1032 470 1151 483
rect 1032 424 1092 470
rect 1138 424 1151 470
rect 1032 411 1151 424
rect 1199 470 1319 483
rect 1199 424 1212 470
rect 1258 424 1319 470
rect 1032 340 1095 411
rect 796 296 916 340
rect 975 296 1095 340
rect 1199 296 1319 424
rect 1467 470 1539 483
rect 1467 424 1480 470
rect 1526 424 1539 470
rect 1467 411 1539 424
rect 1615 470 1715 573
rect 1819 529 1919 573
rect 1615 424 1656 470
rect 1702 424 1715 470
rect 1615 411 1715 424
rect 124 112 244 156
rect 348 112 468 156
rect 572 112 692 156
rect 796 64 916 156
rect 975 112 1095 156
rect 1199 112 1319 156
rect 1467 64 1507 411
rect 1655 321 1715 411
rect 1879 483 1919 529
rect 2257 483 2357 573
rect 2461 529 2561 573
rect 2461 483 2535 529
rect 2665 513 2765 573
rect 2869 513 2969 573
rect 2665 483 2969 513
rect 1879 470 2357 483
rect 1879 424 2052 470
rect 2098 424 2357 470
rect 1879 411 2357 424
rect 1655 277 1775 321
rect 1879 277 1999 411
rect 2247 366 2357 411
rect 2415 470 2535 483
rect 2415 424 2428 470
rect 2474 424 2535 470
rect 2247 322 2367 366
rect 2415 322 2535 424
rect 2639 470 2969 483
rect 2639 424 2652 470
rect 2698 441 2969 470
rect 2698 424 2759 441
rect 2639 322 2759 424
rect 2863 366 2969 441
rect 2863 322 2983 366
rect 1655 93 1775 137
rect 1879 93 1999 137
rect 2247 78 2367 122
rect 2415 78 2535 122
rect 2639 78 2759 122
rect 2863 78 2983 122
rect 796 24 1507 64
<< polycontact >>
rect 142 424 188 470
rect 897 497 943 543
rect 361 424 407 470
rect 689 369 735 415
rect 1092 424 1138 470
rect 1212 424 1258 470
rect 1480 424 1526 470
rect 1656 424 1702 470
rect 2052 424 2098 470
rect 2428 424 2474 470
rect 2652 424 2698 470
<< metal1 >>
rect 0 918 3136 1098
rect 139 839 185 918
rect 139 688 185 699
rect 711 839 757 850
rect 1161 827 1207 918
rect 1744 850 1790 918
rect 1161 770 1207 781
rect 1365 839 1411 850
rect 711 635 757 699
rect 1092 699 1365 724
rect 1744 839 3044 850
rect 1744 827 2590 839
rect 1790 781 2182 827
rect 2228 804 2590 827
rect 1744 770 2228 781
rect 2386 726 2432 737
rect 1411 699 2340 724
rect 1092 678 2340 699
rect 597 589 1046 635
rect 142 470 194 542
rect 188 424 194 470
rect 142 354 194 424
rect 242 424 361 470
rect 407 424 418 470
rect 242 354 418 424
rect 49 261 543 307
rect 49 215 95 261
rect 497 215 543 261
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 597 215 643 589
rect 689 497 897 543
rect 943 497 954 543
rect 689 415 735 497
rect 689 358 735 369
rect 1000 367 1046 589
rect 1092 470 1138 678
rect 1092 413 1138 424
rect 1201 424 1212 470
rect 1258 424 1269 470
rect 1201 367 1269 424
rect 1000 321 1269 367
rect 1124 215 1170 226
rect 597 169 721 215
rect 767 169 778 215
rect 497 158 543 169
rect 1124 90 1170 169
rect 1348 215 1394 678
rect 1480 586 1540 632
rect 1586 586 1597 632
rect 1937 586 1948 632
rect 1994 586 2005 632
rect 1480 470 1526 586
rect 1937 470 1983 586
rect 1645 424 1656 470
rect 1702 424 1983 470
rect 1480 215 1526 424
rect 1804 215 1850 226
rect 1480 169 1580 215
rect 1626 169 1637 215
rect 1348 158 1394 169
rect 1804 90 1850 169
rect 1937 196 1983 424
rect 2046 470 2098 481
rect 2046 424 2052 470
rect 2294 470 2340 678
rect 2636 804 2998 839
rect 2590 688 2636 699
rect 2718 726 2840 737
rect 2432 586 2577 621
rect 2386 575 2577 586
rect 2718 586 2794 726
rect 2998 688 3044 699
rect 2718 578 2840 586
rect 2531 481 2577 575
rect 2531 470 2698 481
rect 2294 424 2428 470
rect 2474 424 2485 470
rect 2531 424 2652 470
rect 2046 242 2098 424
rect 2531 413 2698 424
rect 2531 378 2577 413
rect 2172 332 2577 378
rect 2172 309 2218 332
rect 2788 318 2840 578
rect 1937 150 2028 196
rect 2074 150 2085 196
rect 2718 309 2840 318
rect 2172 158 2218 169
rect 2564 275 2610 286
rect 2718 242 2788 309
rect 2834 169 2840 309
rect 2788 158 2840 169
rect 3012 275 3058 286
rect 2564 90 2610 135
rect 3012 90 3058 135
rect 0 -90 3136 90
<< labels >>
flabel metal1 s 2046 242 2098 481 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel metal1 s 242 354 418 470 0 FreeSans 200 0 0 0 E
port 2 nsew default input
flabel metal1 s 2718 578 2840 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 918 3136 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3012 226 3058 286 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 2788 318 2840 578 1 Q
port 4 nsew default output
rlabel metal1 s 2718 242 2840 318 1 Q
port 4 nsew default output
rlabel metal1 s 2788 158 2840 242 1 Q
port 4 nsew default output
rlabel metal1 s 1744 850 1790 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1161 850 1207 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 139 850 185 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1744 804 3044 850 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1161 804 1207 850 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 139 804 185 850 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2998 770 3044 804 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2590 770 2636 804 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1744 770 2228 804 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1161 770 1207 804 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 139 770 185 804 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2998 688 3044 770 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2590 688 2636 770 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 139 688 185 770 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2564 226 2610 286 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3012 215 3058 226 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2564 215 2610 226 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1804 215 1850 226 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1124 215 1170 226 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3012 90 3058 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2564 90 2610 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1804 90 1850 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1124 90 1170 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 215 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3136 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 1008
string GDS_END 843488
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 836060
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
