magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 4704 844
rect 49 506 95 724
rect 273 611 319 676
rect 466 657 534 724
rect 701 611 747 676
rect 914 657 982 724
rect 1149 611 1195 676
rect 1362 657 1430 724
rect 1597 611 1643 676
rect 1810 657 1878 724
rect 2034 611 2110 676
rect 2258 657 2326 724
rect 2493 611 2539 676
rect 2706 657 2774 724
rect 2941 611 2987 676
rect 3154 657 3222 724
rect 3389 611 3435 676
rect 3602 657 3670 724
rect 3837 611 3883 676
rect 4050 657 4118 724
rect 4285 611 4331 676
rect 273 470 4331 611
rect 4509 506 4555 724
rect 126 348 1980 424
rect 2206 301 2386 470
rect 2504 348 4480 424
rect 262 175 4362 301
rect 49 60 95 140
rect 262 107 330 175
rect 486 60 554 129
rect 710 107 778 175
rect 934 60 1002 129
rect 1158 107 1226 175
rect 1382 60 1450 129
rect 1606 107 1674 175
rect 1830 60 1898 129
rect 2054 107 2122 175
rect 2278 60 2346 129
rect 2502 107 2570 175
rect 2726 60 2794 129
rect 2950 107 3018 175
rect 3174 60 3242 129
rect 3398 107 3466 175
rect 3622 60 3690 129
rect 3846 107 3914 175
rect 4070 60 4138 129
rect 4294 107 4362 175
rect 4518 60 4586 129
rect 0 -60 4704 60
<< labels >>
rlabel metal1 s 126 348 1980 424 6 I
port 1 nsew default input
rlabel metal1 s 2504 348 4480 424 6 I
port 1 nsew default input
rlabel metal1 s 4285 611 4331 676 6 ZN
port 2 nsew default output
rlabel metal1 s 3837 611 3883 676 6 ZN
port 2 nsew default output
rlabel metal1 s 3389 611 3435 676 6 ZN
port 2 nsew default output
rlabel metal1 s 2941 611 2987 676 6 ZN
port 2 nsew default output
rlabel metal1 s 2493 611 2539 676 6 ZN
port 2 nsew default output
rlabel metal1 s 2034 611 2110 676 6 ZN
port 2 nsew default output
rlabel metal1 s 1597 611 1643 676 6 ZN
port 2 nsew default output
rlabel metal1 s 1149 611 1195 676 6 ZN
port 2 nsew default output
rlabel metal1 s 701 611 747 676 6 ZN
port 2 nsew default output
rlabel metal1 s 273 611 319 676 6 ZN
port 2 nsew default output
rlabel metal1 s 273 470 4331 611 6 ZN
port 2 nsew default output
rlabel metal1 s 2206 301 2386 470 6 ZN
port 2 nsew default output
rlabel metal1 s 262 175 4362 301 6 ZN
port 2 nsew default output
rlabel metal1 s 4294 107 4362 175 6 ZN
port 2 nsew default output
rlabel metal1 s 3846 107 3914 175 6 ZN
port 2 nsew default output
rlabel metal1 s 3398 107 3466 175 6 ZN
port 2 nsew default output
rlabel metal1 s 2950 107 3018 175 6 ZN
port 2 nsew default output
rlabel metal1 s 2502 107 2570 175 6 ZN
port 2 nsew default output
rlabel metal1 s 2054 107 2122 175 6 ZN
port 2 nsew default output
rlabel metal1 s 1606 107 1674 175 6 ZN
port 2 nsew default output
rlabel metal1 s 1158 107 1226 175 6 ZN
port 2 nsew default output
rlabel metal1 s 710 107 778 175 6 ZN
port 2 nsew default output
rlabel metal1 s 262 107 330 175 6 ZN
port 2 nsew default output
rlabel metal1 s 0 724 4704 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 657 4555 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4050 657 4118 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3602 657 3670 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3154 657 3222 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2706 657 2774 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2258 657 2326 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1810 657 1878 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1362 657 1430 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 914 657 982 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 466 657 534 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 657 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 506 4555 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 129 95 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4518 60 4586 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 129 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4704 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4704 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 840698
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 830502
<< end >>
