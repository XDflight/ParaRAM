magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 2209 5116 4648 6727
rect 2137 5115 4648 5116
rect 2101 4660 4696 5115
<< psubdiff >>
rect 1993 6997 5034 7162
rect 1835 2102 1995 2103
rect 1835 2043 2627 2102
rect 1835 1997 1892 2043
rect 1938 1997 2050 2043
rect 2096 1997 2208 2043
rect 2254 1997 2366 2043
rect 2412 1997 2524 2043
rect 2570 1997 2627 2043
rect 1835 1937 2627 1997
rect 2468 1756 2627 1937
rect 4875 1055 5034 6997
rect 4875 1009 4932 1055
rect 4978 1009 5034 1055
rect 4875 892 5034 1009
rect 4875 846 4932 892
rect 4978 846 5034 892
rect 4875 728 5034 846
rect 4875 682 4932 728
rect 4978 682 5034 728
rect 4875 565 5034 682
rect 4875 519 4932 565
rect 4978 519 5034 565
rect 2468 235 2627 416
rect 4875 402 5034 519
rect 4875 356 4932 402
rect 4978 356 5034 402
rect 2468 234 2628 235
rect 4875 234 5034 356
rect 2468 69 5034 234
<< nsubdiff >>
rect 2245 4911 2400 4968
rect 2245 4865 2299 4911
rect 2345 4865 2400 4911
rect 2245 4808 2400 4865
rect 4398 4911 4553 4968
rect 4398 4865 4452 4911
rect 4498 4865 4553 4911
rect 4398 4808 4553 4865
<< psubdiffcont >>
rect 1892 1997 1938 2043
rect 2050 1997 2096 2043
rect 2208 1997 2254 2043
rect 2366 1997 2412 2043
rect 2524 1997 2570 2043
rect 4932 1009 4978 1055
rect 4932 846 4978 892
rect 4932 682 4978 728
rect 4932 519 4978 565
rect 4932 356 4978 402
<< nsubdiffcont >>
rect 2299 4865 2345 4911
rect 4452 4865 4498 4911
<< polysilicon >>
rect 3151 6740 3719 6759
rect 3151 6694 3412 6740
rect 3458 6694 3719 6740
rect 3151 6659 3719 6694
rect 2464 5746 2584 6106
rect 2688 5746 2808 6106
rect 3375 5746 3494 6061
rect 4049 5746 4169 6106
rect 4273 5746 4393 6106
rect 2095 5216 2179 5235
rect 2095 5170 2114 5216
rect 2160 5206 2179 5216
rect 4635 5216 4719 5235
rect 4049 5206 4169 5207
rect 4273 5206 4393 5207
rect 4635 5206 4654 5216
rect 2160 5170 2808 5206
rect 2095 5151 2808 5170
rect 4049 5170 4654 5206
rect 4700 5170 4719 5216
rect 4049 5151 4719 5170
rect 2699 4721 2917 4740
rect 2699 4675 2718 4721
rect 2764 4675 2917 4721
rect 2699 4656 2917 4675
rect 3021 4621 3141 4738
rect 2556 4507 2760 4526
rect 2556 4461 2695 4507
rect 2741 4461 2760 4507
rect 2556 4442 2760 4461
rect 2556 3950 2676 4442
rect 3021 4310 3124 4621
rect 3245 4507 3365 4818
rect 3245 4461 3264 4507
rect 3310 4461 3365 4507
rect 3021 4291 3159 4310
rect 3021 4267 3094 4291
rect 2780 4245 3094 4267
rect 3140 4245 3159 4291
rect 2780 4226 3159 4245
rect 2780 4197 3124 4226
rect 2780 3950 2900 4197
rect 3004 3953 3124 4197
rect 3245 4105 3365 4461
rect 3487 4619 3589 4769
rect 3720 4623 3813 4818
rect 3917 4723 4121 4742
rect 3917 4677 4056 4723
rect 4102 4677 4121 4723
rect 3917 4658 4121 4677
rect 3487 4507 3615 4619
rect 3487 4461 3550 4507
rect 3596 4461 3615 4507
rect 3487 4108 3615 4461
rect 3720 4291 3848 4623
rect 3720 4245 3739 4291
rect 3785 4267 3848 4291
rect 4124 4507 4244 4526
rect 4124 4461 4143 4507
rect 4189 4461 4244 4507
rect 3785 4245 4020 4267
rect 3720 4197 4020 4245
rect 3245 3989 3348 4105
rect 3487 3950 3572 4108
rect 3720 4101 3848 4197
rect 3720 3957 3796 4101
rect 3900 3950 4020 4197
rect 4124 3957 4244 4461
rect 2257 3208 2450 3253
rect 2257 3162 2331 3208
rect 2377 3162 2450 3208
rect 2257 3116 2450 3162
rect 4418 3208 4611 3253
rect 4418 3162 4492 3208
rect 4538 3162 4611 3208
rect 4418 3116 4611 3162
rect 2589 2401 4277 2447
rect 2589 2355 2663 2401
rect 2709 2355 2966 2401
rect 3012 2355 3412 2401
rect 3458 2355 3864 2401
rect 3910 2355 4156 2401
rect 4202 2355 4277 2401
rect 2589 2309 4277 2355
rect 3034 1595 3154 1708
rect 3034 1593 3378 1595
rect 2870 1574 3378 1593
rect 2870 1528 2889 1574
rect 3029 1534 3378 1574
rect 3029 1528 3154 1534
rect 2870 1509 3154 1528
rect 3034 1382 3154 1509
rect 3258 1352 3378 1534
rect 3482 1593 3602 1672
rect 3706 1642 3826 1672
rect 3706 1593 4050 1642
rect 3482 1588 4050 1593
rect 3482 1574 3826 1588
rect 3482 1528 3549 1574
rect 3689 1528 3826 1574
rect 3482 1509 3826 1528
rect 3482 1387 3602 1509
rect 3706 1378 3826 1509
rect 4154 1581 4274 1640
rect 4154 1562 4449 1581
rect 4154 1516 4290 1562
rect 4430 1516 4449 1562
rect 4154 1497 4449 1516
rect 4154 1452 4274 1497
rect 3930 1391 4274 1452
rect 3930 1353 4050 1391
rect 4154 1378 4274 1391
<< polycontact >>
rect 3412 6694 3458 6740
rect 2114 5170 2160 5216
rect 4654 5170 4700 5216
rect 2718 4675 2764 4721
rect 2695 4461 2741 4507
rect 3264 4461 3310 4507
rect 3094 4245 3140 4291
rect 4056 4677 4102 4723
rect 3550 4461 3596 4507
rect 3739 4245 3785 4291
rect 4143 4461 4189 4507
rect 2331 3162 2377 3208
rect 4492 3162 4538 3208
rect 2663 2355 2709 2401
rect 2966 2355 3012 2401
rect 3412 2355 3458 2401
rect 3864 2355 3910 2401
rect 4156 2355 4202 2401
rect 2889 1528 3029 1574
rect 3549 1528 3689 1574
rect 4290 1516 4430 1562
<< metal1 >>
rect 1756 8029 2524 8033
rect 1756 8009 2633 8029
rect 1756 7957 2355 8009
rect 2407 7957 2541 8009
rect 2593 7957 2633 8009
rect 1756 7937 2633 7957
rect 3076 8009 4501 8033
rect 3076 7957 4219 8009
rect 4271 7957 4405 8009
rect 4457 7957 4501 8009
rect 1756 7936 2524 7937
rect 3076 7936 4501 7957
rect 2430 7824 2524 7936
rect 2430 7800 4501 7824
rect 2430 7748 2737 7800
rect 2789 7748 2923 7800
rect 2975 7748 3541 7800
rect 3593 7748 3727 7800
rect 3779 7748 4501 7800
rect 2430 7727 4501 7748
rect 1756 7478 4885 7616
rect 1251 7339 4501 7362
rect 1251 7287 3410 7339
rect 3462 7287 4501 7339
rect 1251 7265 4501 7287
rect 1844 7006 5025 7153
rect 3271 6823 3609 6899
rect 3387 6822 3482 6823
rect 2797 6741 2925 6763
rect 3388 6750 3482 6822
rect 1844 2094 1986 6741
rect 2387 6740 3310 6741
rect 2387 6688 2835 6740
rect 2887 6688 3310 6740
rect 2387 6666 3310 6688
rect 2387 6577 2458 6666
rect 2386 6132 2458 6577
rect 2596 6424 2688 6464
rect 2596 6372 2616 6424
rect 2668 6372 2688 6424
rect 2596 6238 2688 6372
rect 2596 6186 2616 6238
rect 2668 6186 2688 6238
rect 2596 6145 2688 6186
rect 2837 6132 2883 6666
rect 3239 6464 3310 6666
rect 3388 6698 3408 6750
rect 3460 6698 3482 6750
rect 3388 6694 3412 6698
rect 3458 6694 3482 6698
rect 3388 6657 3482 6694
rect 3559 6718 4483 6741
rect 3559 6666 3970 6718
rect 4022 6666 4483 6718
rect 3559 6464 3631 6666
rect 3932 6644 4060 6666
rect 3239 6424 3369 6464
rect 3239 6372 3297 6424
rect 3349 6372 3369 6424
rect 3239 6238 3369 6372
rect 3239 6186 3297 6238
rect 3349 6186 3369 6238
rect 3239 6145 3369 6186
rect 3503 6424 3631 6464
rect 3503 6372 3523 6424
rect 3575 6372 3631 6424
rect 3503 6238 3631 6372
rect 3503 6186 3523 6238
rect 3575 6186 3631 6238
rect 3503 6145 3631 6186
rect 3239 6140 3310 6145
rect 3559 6140 3631 6145
rect 3939 6140 4055 6644
rect 4181 6424 4273 6464
rect 4181 6372 4201 6424
rect 4253 6372 4273 6424
rect 4181 6238 4273 6372
rect 4181 6186 4201 6238
rect 4253 6186 4273 6238
rect 4181 6145 4273 6186
rect 4411 6140 4483 6666
rect 2378 5884 2467 6061
rect 2843 5884 2933 6061
rect 3278 6057 4468 6061
rect 3276 6036 4468 6057
rect 3276 5984 3316 6036
rect 3368 5984 4468 6036
rect 3276 5968 4468 5984
rect 3276 5964 3404 5968
rect 3467 5884 3595 5885
rect 2378 5864 3595 5884
rect 2378 5812 3503 5864
rect 3555 5812 3595 5864
rect 2378 5792 3595 5812
rect 2378 5791 3591 5792
rect 2378 5711 2467 5791
rect 2377 5304 2467 5711
rect 2064 5216 2171 5227
rect 2064 5170 2114 5216
rect 2160 5170 2171 5216
rect 2613 5195 2659 5349
rect 2837 5266 2883 5791
rect 3974 5370 4020 5968
rect 3300 5195 3346 5349
rect 2064 5159 2171 5170
rect 2064 2438 2136 5159
rect 2448 5120 3346 5195
rect 3524 5195 3570 5274
rect 4198 5195 4244 5349
rect 4422 5304 4468 5968
rect 4643 5216 4916 5227
rect 3524 5120 4340 5195
rect 4643 5170 4654 5216
rect 4700 5170 4916 5216
rect 4643 5159 4916 5170
rect 2286 5024 2380 5025
rect 2264 4911 2380 5024
rect 2264 4865 2299 4911
rect 2345 4865 2380 4911
rect 2264 4719 2380 4865
rect 2448 4319 2520 5120
rect 3151 5024 3245 5025
rect 3623 5024 3717 5025
rect 2679 4721 2794 4975
rect 2679 4675 2718 4721
rect 2764 4675 2794 4721
rect 2679 4664 2794 4675
rect 2911 4532 2975 4984
rect 3144 4719 3260 5024
rect 3398 4809 3471 4975
rect 2684 4510 2992 4532
rect 2684 4507 2722 4510
rect 2684 4461 2695 4507
rect 2684 4458 2722 4461
rect 2774 4458 2902 4510
rect 2954 4458 2992 4510
rect 2684 4436 2992 4458
rect 3083 4510 3329 4544
rect 3083 4458 3231 4510
rect 3283 4507 3329 4510
rect 3310 4461 3329 4507
rect 3283 4458 3329 4461
rect 2332 4298 2520 4319
rect 2332 4246 2428 4298
rect 2480 4246 2520 4298
rect 2332 4226 2520 4246
rect 2332 4145 2403 4226
rect 2332 4071 2518 4145
rect 2213 3244 2329 3988
rect 2446 3910 2518 4071
rect 2911 3891 2975 4436
rect 3083 4424 3329 4458
rect 3083 4299 3293 4326
rect 3399 4322 3471 4809
rect 3610 4719 3725 5024
rect 3539 4510 3758 4544
rect 3886 4532 3958 4973
rect 4039 4723 4155 4984
rect 4039 4677 4056 4723
rect 4102 4677 4155 4723
rect 4039 4664 4155 4677
rect 3539 4507 3587 4510
rect 3539 4461 3550 4507
rect 3539 4458 3587 4461
rect 3639 4458 3758 4510
rect 3539 4424 3758 4458
rect 3883 4510 4200 4532
rect 3883 4458 3921 4510
rect 3973 4458 4101 4510
rect 4153 4507 4200 4510
rect 4189 4461 4200 4507
rect 4153 4458 4200 4461
rect 3883 4436 4200 4458
rect 4268 4530 4340 5120
rect 4418 5024 4512 5025
rect 4418 4911 4534 5024
rect 4418 4865 4452 4911
rect 4498 4865 4534 4911
rect 4418 4719 4534 4865
rect 4268 4509 4396 4530
rect 4268 4457 4304 4509
rect 4356 4457 4396 4509
rect 4268 4437 4396 4457
rect 3083 4291 3121 4299
rect 3083 4245 3094 4291
rect 3173 4247 3293 4299
rect 3140 4245 3293 4247
rect 3083 4202 3293 4245
rect 3371 4299 3499 4322
rect 3371 4247 3409 4299
rect 3461 4247 3499 4299
rect 3371 4225 3499 4247
rect 3577 4299 3796 4326
rect 3577 4247 3697 4299
rect 3749 4291 3796 4299
rect 3577 4245 3739 4247
rect 3785 4245 3796 4291
rect 3399 3988 3471 4225
rect 3577 4202 3796 4245
rect 3886 3999 3958 4436
rect 4268 4227 4340 4437
rect 4475 4322 4547 4533
rect 4474 4319 4547 4322
rect 4440 4298 4568 4319
rect 4440 4246 4476 4298
rect 4528 4246 4568 4298
rect 4440 4226 4568 4246
rect 4474 4225 4547 4226
rect 4475 4145 4547 4225
rect 3398 3855 3471 3988
rect 3826 3891 3958 3999
rect 4273 4071 4547 4145
rect 4273 3910 4319 4071
rect 2679 3245 2794 3411
rect 3144 3245 3260 3411
rect 3610 3245 3725 3411
rect 4075 3410 4095 3411
rect 4049 3245 4095 3410
rect 4541 3245 4657 3988
rect 2213 3242 2411 3244
rect 2213 3221 2486 3242
rect 2213 3208 2394 3221
rect 2213 3162 2331 3208
rect 2377 3169 2394 3208
rect 2446 3169 2486 3221
rect 2377 3162 2486 3169
rect 2213 3149 2486 3162
rect 2679 3152 4095 3245
rect 4540 3244 4657 3245
rect 4457 3242 4657 3244
rect 4378 3221 4657 3242
rect 4378 3169 4414 3221
rect 4466 3208 4657 3221
rect 4466 3169 4492 3208
rect 4378 3162 4492 3169
rect 4538 3162 4657 3208
rect 2213 3125 2411 3149
rect 2703 2518 2818 3152
rect 3151 2518 3266 3152
rect 3599 2518 3714 3152
rect 4047 2518 4162 3152
rect 4378 3149 4657 3162
rect 4457 3125 4657 3149
rect 4844 2438 4916 5159
rect 2064 2401 4916 2438
rect 2064 2355 2663 2401
rect 2709 2355 2966 2401
rect 3012 2355 3412 2401
rect 3458 2355 3864 2401
rect 3910 2355 4156 2401
rect 4202 2355 4916 2401
rect 2064 2318 4916 2355
rect 1844 2093 1987 2094
rect 1844 2043 2619 2093
rect 1844 1997 1892 2043
rect 1938 1997 2050 2043
rect 2096 1997 2208 2043
rect 2254 1997 2366 2043
rect 2412 1997 2524 2043
rect 2570 1997 2619 2043
rect 1844 1946 2619 1997
rect 2477 225 2619 1946
rect 3386 1990 3478 2030
rect 3386 1938 3406 1990
rect 3458 1938 3478 1990
rect 3386 1804 3478 1938
rect 2749 1577 3057 1597
rect 2749 1525 2779 1577
rect 2831 1574 2965 1577
rect 3017 1574 3057 1577
rect 2831 1528 2889 1574
rect 3029 1528 3057 1574
rect 2831 1525 2965 1528
rect 3017 1525 3057 1528
rect 2749 1505 3057 1525
rect 3183 1585 3229 1762
rect 3386 1752 3406 1804
rect 3458 1752 3478 1804
rect 3386 1711 3478 1752
rect 3828 1990 3920 2030
rect 3828 1938 3848 1990
rect 3900 1938 3920 1990
rect 3828 1804 3920 1938
rect 3828 1752 3848 1804
rect 3900 1752 3920 1804
rect 3828 1711 3920 1752
rect 4276 1990 4368 2030
rect 4276 1938 4296 1990
rect 4348 1938 4368 1990
rect 4276 1804 4368 1938
rect 4276 1752 4296 1804
rect 4348 1752 4368 1804
rect 4276 1711 4368 1752
rect 3183 1574 3700 1585
rect 3183 1528 3549 1574
rect 3689 1528 3700 1574
rect 3183 1517 3700 1528
rect 4251 1566 4559 1586
rect 2925 545 3040 1331
rect 3183 1293 3229 1517
rect 4251 1514 4281 1566
rect 4333 1562 4467 1566
rect 4430 1516 4467 1562
rect 4333 1514 4467 1516
rect 4519 1514 4559 1566
rect 4251 1494 4559 1514
rect 3373 661 3488 1331
rect 3601 1296 3693 1336
rect 3601 1244 3621 1296
rect 3673 1244 3693 1296
rect 3601 1110 3693 1244
rect 3601 1058 3621 1110
rect 3673 1058 3693 1110
rect 3601 1017 3693 1058
rect 2924 541 3040 545
rect 3372 541 3488 661
rect 3820 541 3936 1331
rect 4061 1296 4153 1336
rect 4061 1244 4081 1296
rect 4133 1244 4153 1296
rect 4061 1110 4153 1244
rect 4061 1058 4081 1110
rect 4133 1058 4153 1110
rect 4061 1017 4153 1058
rect 4268 541 4384 1331
rect 4883 1055 5025 1155
rect 4883 1009 4932 1055
rect 4978 1009 5025 1055
rect 4883 892 5025 1009
rect 4883 846 4932 892
rect 4978 846 5025 892
rect 4883 728 5025 846
rect 4883 682 4932 728
rect 4978 682 5025 728
rect 4883 565 5025 682
rect 4883 519 4932 565
rect 4978 519 5025 565
rect 4883 402 5025 519
rect 4883 356 4932 402
rect 4978 356 5025 402
rect 4883 225 5025 356
rect 2477 78 5025 225
<< via1 >>
rect 2355 7957 2407 8009
rect 2541 7957 2593 8009
rect 4219 7957 4271 8009
rect 4405 7957 4457 8009
rect 2737 7748 2789 7800
rect 2923 7748 2975 7800
rect 3541 7748 3593 7800
rect 3727 7748 3779 7800
rect 3410 7287 3462 7339
rect 2835 6688 2887 6740
rect 2616 6372 2668 6424
rect 2616 6186 2668 6238
rect 3408 6740 3460 6750
rect 3408 6698 3412 6740
rect 3412 6698 3458 6740
rect 3458 6698 3460 6740
rect 3970 6666 4022 6718
rect 3297 6372 3349 6424
rect 3297 6186 3349 6238
rect 3523 6372 3575 6424
rect 3523 6186 3575 6238
rect 4201 6372 4253 6424
rect 4201 6186 4253 6238
rect 3316 5984 3368 6036
rect 3503 5812 3555 5864
rect 2722 4507 2774 4510
rect 2722 4461 2741 4507
rect 2741 4461 2774 4507
rect 2722 4458 2774 4461
rect 2902 4458 2954 4510
rect 3231 4507 3283 4510
rect 3231 4461 3264 4507
rect 3264 4461 3283 4507
rect 3231 4458 3283 4461
rect 2428 4246 2480 4298
rect 3587 4507 3639 4510
rect 3587 4461 3596 4507
rect 3596 4461 3639 4507
rect 3587 4458 3639 4461
rect 3921 4458 3973 4510
rect 4101 4507 4153 4510
rect 4101 4461 4143 4507
rect 4143 4461 4153 4507
rect 4101 4458 4153 4461
rect 4304 4457 4356 4509
rect 3121 4291 3173 4299
rect 3121 4247 3140 4291
rect 3140 4247 3173 4291
rect 3409 4247 3461 4299
rect 3697 4291 3749 4299
rect 3697 4247 3739 4291
rect 3739 4247 3749 4291
rect 4476 4246 4528 4298
rect 2394 3169 2446 3221
rect 4414 3169 4466 3221
rect 3406 1938 3458 1990
rect 2779 1525 2831 1577
rect 2965 1574 3017 1577
rect 2965 1528 3017 1574
rect 2965 1525 3017 1528
rect 3406 1752 3458 1804
rect 3848 1938 3900 1990
rect 3848 1752 3900 1804
rect 4296 1938 4348 1990
rect 4296 1752 4348 1804
rect 4281 1562 4333 1566
rect 4281 1516 4290 1562
rect 4290 1516 4333 1562
rect 4281 1514 4333 1516
rect 4467 1514 4519 1566
rect 3621 1244 3673 1296
rect 3621 1058 3673 1110
rect 4081 1244 4133 1296
rect 4081 1058 4133 1110
<< metal2 >>
rect 2433 8033 2522 8146
rect 3052 8033 3141 8146
rect 2432 8029 2522 8033
rect 2325 8009 2633 8029
rect 2325 7957 2355 8009
rect 2407 7957 2541 8009
rect 2593 7957 2633 8009
rect 2325 7937 2633 7957
rect 2432 7936 2522 7937
rect 3051 7936 3141 8033
rect 2812 7820 2906 7824
rect 3671 7820 3761 8146
rect 4290 8033 4380 8146
rect 3950 8029 4380 8033
rect 3950 8009 4497 8029
rect 3950 7957 4219 8009
rect 4271 7957 4405 8009
rect 4457 7957 4497 8009
rect 3950 7937 4497 7957
rect 3950 7936 4380 7937
rect 1684 7802 1992 7820
rect 1684 7746 1712 7802
rect 1768 7746 1898 7802
rect 1954 7746 1992 7802
rect 1684 7728 1992 7746
rect 2707 7800 3015 7820
rect 2707 7748 2737 7800
rect 2789 7748 2923 7800
rect 2975 7748 3015 7800
rect 2707 7728 3015 7748
rect 3511 7800 3819 7820
rect 3511 7748 3541 7800
rect 3593 7748 3727 7800
rect 3779 7748 3819 7800
rect 3511 7728 3819 7748
rect 2812 7727 2906 7728
rect 3671 7727 3761 7728
rect 2813 6763 2906 7727
rect 3373 7339 3501 7362
rect 3373 7287 3410 7339
rect 3462 7287 3501 7339
rect 3373 7265 3501 7287
rect 2798 6740 2926 6763
rect 2798 6688 2835 6740
rect 2887 6688 2926 6740
rect 2798 6666 2926 6688
rect 3388 6750 3482 7265
rect 3388 6698 3408 6750
rect 3460 6698 3482 6750
rect 3950 6741 4044 7936
rect 3388 6657 3482 6698
rect 3933 6718 4061 6741
rect 3933 6666 3970 6718
rect 4022 6666 4061 6718
rect 3933 6644 4061 6666
rect 2595 6424 2688 6464
rect 2595 6372 2616 6424
rect 2668 6372 2688 6424
rect 2595 6238 2688 6372
rect 2595 6186 2616 6238
rect 2668 6186 2688 6238
rect 2595 6146 2688 6186
rect 3277 6424 3369 6464
rect 3277 6372 3297 6424
rect 3349 6372 3369 6424
rect 3277 6238 3369 6372
rect 3277 6186 3297 6238
rect 3349 6186 3369 6238
rect 3277 6172 3369 6186
rect 3503 6424 3595 6464
rect 3503 6372 3523 6424
rect 3575 6372 3595 6424
rect 3503 6238 3595 6372
rect 3503 6186 3523 6238
rect 3575 6186 3595 6238
rect 3503 6172 3595 6186
rect 4181 6424 4274 6464
rect 4181 6372 4201 6424
rect 4253 6372 4274 6424
rect 4181 6238 4274 6372
rect 4181 6186 4201 6238
rect 4253 6186 4274 6238
rect 2595 6061 2685 6146
rect 2071 5968 2685 6061
rect 3276 6057 3370 6172
rect 3276 6036 3403 6057
rect 3276 5984 3316 6036
rect 3368 5984 3403 6036
rect 2071 4533 2160 5968
rect 3276 5964 3403 5984
rect 3276 5791 3370 5964
rect 3502 5885 3596 6172
rect 4181 6063 4274 6186
rect 4181 5966 4696 6063
rect 3468 5864 3596 5885
rect 3468 5812 3503 5864
rect 3555 5812 3596 5864
rect 3468 5792 3596 5812
rect 3502 5791 3596 5792
rect 2071 4510 4461 4533
rect 2071 4458 2722 4510
rect 2774 4458 2902 4510
rect 2954 4458 3231 4510
rect 3283 4458 3587 4510
rect 3639 4458 3921 4510
rect 3973 4458 4101 4510
rect 4153 4509 4461 4510
rect 4153 4458 4304 4509
rect 2071 4457 4304 4458
rect 4356 4457 4461 4509
rect 2071 4436 4461 4457
rect 2071 2309 2160 4436
rect 4602 4322 4696 5966
rect 2388 4299 4696 4322
rect 2388 4298 3121 4299
rect 2388 4246 2428 4298
rect 2480 4247 3121 4298
rect 3173 4247 3409 4299
rect 3461 4247 3697 4299
rect 3749 4298 4696 4299
rect 3749 4247 4476 4298
rect 2480 4246 4476 4247
rect 4528 4246 4696 4298
rect 2388 4225 4696 4246
rect 2358 3221 2698 3245
rect 2358 3150 2394 3221
rect 2446 3206 2698 3221
rect 2450 3150 2606 3206
rect 2662 3150 2698 3206
rect 2358 3111 2698 3150
rect 4167 3221 4507 3245
rect 4167 3206 4414 3221
rect 4466 3206 4507 3221
rect 4167 3150 4203 3206
rect 4259 3169 4414 3206
rect 4259 3150 4415 3169
rect 4471 3150 4507 3206
rect 4167 3111 4507 3150
rect 4602 2311 4696 4225
rect 2071 2216 2838 2309
rect 2749 1597 2838 2216
rect 4279 2214 4907 2311
rect 3386 1990 3479 2030
rect 3386 1938 3406 1990
rect 3458 1938 3479 1990
rect 3386 1804 3479 1938
rect 3386 1752 3406 1804
rect 3458 1781 3479 1804
rect 3827 1990 3921 2030
rect 3827 1938 3848 1990
rect 3900 1938 3921 1990
rect 3827 1804 3921 1938
rect 3458 1780 3480 1781
rect 3827 1780 3848 1804
rect 3458 1752 3848 1780
rect 3900 1752 3921 1804
rect 4275 1990 4369 2030
rect 4275 1938 4296 1990
rect 4348 1938 4369 1990
rect 4275 1804 4369 1938
rect 4275 1780 4296 1804
rect 3386 1683 3921 1752
rect 4060 1752 4296 1780
rect 4348 1752 4369 1804
rect 4060 1683 4369 1752
rect 2749 1577 3057 1597
rect 2749 1525 2779 1577
rect 2831 1525 2965 1577
rect 3017 1525 3057 1577
rect 2749 1505 3057 1525
rect 2749 1504 2838 1505
rect 3601 1296 3695 1683
rect 3601 1244 3621 1296
rect 3673 1244 3695 1296
rect 3601 1110 3695 1244
rect 3601 1058 3621 1110
rect 3673 1058 3695 1110
rect 3601 -196 3695 1058
rect 4060 1296 4154 1683
rect 4466 1586 4560 2214
rect 4251 1566 4560 1586
rect 4251 1514 4281 1566
rect 4333 1514 4467 1566
rect 4519 1514 4560 1566
rect 4251 1504 4560 1514
rect 4251 1494 4559 1504
rect 4060 1244 4081 1296
rect 4133 1244 4154 1296
rect 4060 1110 4154 1244
rect 4060 1058 4081 1110
rect 4133 1058 4154 1110
rect 4060 -196 4154 1058
<< via2 >>
rect 1712 7746 1768 7802
rect 1898 7746 1954 7802
rect 2394 3169 2446 3206
rect 2446 3169 2450 3206
rect 2394 3150 2450 3169
rect 2606 3150 2662 3206
rect 4203 3150 4259 3206
rect 4415 3169 4466 3206
rect 4466 3169 4471 3206
rect 4415 3150 4471 3169
<< metal3 >>
rect 2430 7936 3130 8033
rect 2430 7824 2524 7936
rect 1684 7802 2524 7824
rect 1684 7746 1712 7802
rect 1768 7746 1898 7802
rect 1954 7746 2524 7802
rect 1684 7727 2524 7746
rect -356 4383 4955 7106
rect -356 3206 5006 4097
rect -356 3150 2394 3206
rect 2450 3150 2606 3206
rect 2662 3150 4203 3206
rect 4259 3150 4415 3206
rect 4471 3150 5006 3206
rect -356 951 5006 3150
rect -357 817 5006 951
rect -356 695 5006 817
rect -356 -172 5006 545
use M1_NWELL06_512x8m81  M1_NWELL06_512x8m81_0
timestamp 1666464484
transform 1 0 3667 0 1 601
box -853 -228 853 228
use M1_NWELL_01_R90_512x8m81  M1_NWELL_01_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 2322 1 0 4888
box 0 0 1 1
use M1_NWELL_01_R90_512x8m81  M1_NWELL_01_R90_512x8m81_1
timestamp 1666464484
transform 0 -1 4475 1 0 4888
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_0
timestamp 1666464484
transform -1 0 3887 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_1
timestamp 1666464484
transform -1 0 4179 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_2
timestamp 1666464484
transform 1 0 4515 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_3
timestamp 1666464484
transform -1 0 2989 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_4
timestamp 1666464484
transform 1 0 2354 0 1 3185
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_5
timestamp 1666464484
transform 1 0 2686 0 1 2378
box 0 0 1 1
use M1_POLY2$$44753964_512x8m81  M1_POLY2$$44753964_512x8m81_6
timestamp 1666464484
transform -1 0 3435 0 1 2378
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1666464484
transform 1 0 3287 0 1 4484
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1666464484
transform 1 0 3117 0 1 4268
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1666464484
transform 1 0 2741 0 1 4698
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1666464484
transform 1 0 2137 0 1 5193
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1666464484
transform 1 0 2718 0 1 4484
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1666464484
transform 1 0 3762 0 1 4268
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1666464484
transform 1 0 3573 0 1 4484
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1666464484
transform 1 0 4166 0 1 4484
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_8
timestamp 1666464484
transform 1 0 4079 0 1 4700
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_9
timestamp 1666464484
transform 1 0 4677 0 1 5193
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_10
timestamp 1666464484
transform 1 0 3435 0 1 6717
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1666464484
transform 1 0 3619 0 1 1551
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1666464484
transform 1 0 4360 0 1 1539
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1666464484
transform 1 0 2959 0 1 1551
box 0 0 1 1
use M1_PSUB$$46555180_512x8m81  M1_PSUB$$46555180_512x8m81_0
timestamp 1666464484
transform 1 0 3439 0 1 7080
box -1424 -83 1424 82
use M1_PSUB$$46556204_512x8m81  M1_PSUB$$46556204_512x8m81_0
timestamp 1666464484
transform 1 0 1915 0 1 4550
box -80 -2613 80 2612
use M1_PSUB$$46557228_512x8m81  M1_PSUB$$46557228_512x8m81_0
timestamp 1666464484
transform 1 0 2231 0 1 2020
box 0 0 1 1
use M1_PSUB$$46558252_512x8m81  M1_PSUB$$46558252_512x8m81_0
timestamp 1666464484
transform 1 0 3674 0 1 152
box -950 -83 950 82
use M1_PSUB_04_R90_512x8m81  M1_PSUB_04_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 2547 1 0 1031
box -817 -80 817 79
use M3_M2$$43371564_512x8m81  M3_M2$$43371564_512x8m81_0
timestamp 1666464484
transform 1 0 4337 0 1 3178
box 0 0 1 1
use M3_M2$$43371564_512x8m81  M3_M2$$43371564_512x8m81_1
timestamp 1666464484
transform 1 0 2528 0 1 3178
box 0 0 1 1
use nmos_1p2$$45107244_512x8m81  nmos_1p2$$45107244_512x8m81_0
timestamp 1666464484
transform -1 0 4243 0 -1 2156
box -119 -73 849 526
use nmos_1p2$$46550060_512x8m81  nmos_1p2$$46550060_512x8m81_0
timestamp 1666464484
transform 1 0 2620 0 1 2510
box -119 -74 1745 640
use nmos_1p2$$46551084_512x8m81  nmos_1p2$$46551084_512x8m81_0
timestamp 1666464484
transform -1 0 3123 0 -1 2156
box -119 -73 177 527
use nmos_1p2$$46552108_512x8m81  nmos_1p2$$46552108_512x8m81_0
timestamp 1666464484
transform 1 0 2587 0 1 3317
box -119 -74 1745 754
use nmos_1p2$$46553132_512x8m81  nmos_1p2$$46553132_512x8m81_0
timestamp 1666464484
transform 1 0 4379 0 1 3317
box -119 -74 177 753
use nmos_1p2$$46553132_512x8m81  nmos_1p2$$46553132_512x8m81_1
timestamp 1666464484
transform 1 0 2363 0 1 3317
box -119 -74 177 753
use pmos_1p2$$46285868_512x8m81  pmos_1p2$$46285868_512x8m81_0
timestamp 1666464484
transform 1 0 3406 0 1 5266
box -286 -142 344 595
use pmos_1p2$$46286892_512x8m81  pmos_1p2$$46286892_512x8m81_0
timestamp 1666464484
transform 1 0 3182 0 1 6132
box -286 -142 792 595
use pmos_1p2$$46549036_512x8m81  pmos_1p2$$46549036_512x8m81_0
timestamp 1666464484
transform -1 0 4243 0 -1 1331
box -286 -142 1463 595
use pmos_1p2$$46896172_512x8m81  pmos_1p2$$46896172_512x8m81_0
timestamp 1666464484
transform 1 0 3052 0 1 4802
box -286 -142 1051 323
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_0
timestamp 1666464484
transform 1 0 2495 0 1 6132
box -286 -142 568 595
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_1
timestamp 1666464484
transform 1 0 2495 0 1 5266
box -286 -142 568 595
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_2
timestamp 1666464484
transform 1 0 4080 0 1 6132
box -286 -142 568 595
use pmos_1p2$$46897196_512x8m81  pmos_1p2$$46897196_512x8m81_3
timestamp 1666464484
transform 1 0 4080 0 1 5266
box -286 -142 568 595
use pmos_1p2$$46898220_512x8m81  pmos_1p2$$46898220_512x8m81_0
timestamp 1666464484
transform 1 0 2828 0 1 4802
box -286 -142 352 323
use pmos_1p2$$46898220_512x8m81  pmos_1p2$$46898220_512x8m81_1
timestamp 1666464484
transform 1 0 3948 0 1 4802
box -286 -142 352 323
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1666464484
transform 1 0 4909 0 1 827
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1666464484
transform 1 0 3834 0 1 2621
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1666464484
transform -1 0 3700 0 -1 2201
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1666464484
transform -1 0 4146 0 -1 2201
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1666464484
transform 1 0 4271 0 1 2621
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1666464484
transform 1 0 3386 0 1 2621
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1666464484
transform -1 0 3033 0 -1 2029
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1666464484
transform 1 0 2523 0 1 827
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1666464484
transform 1 0 2523 0 1 1630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1666464484
transform 1 0 2501 0 1 2621
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1666464484
transform 1 0 2938 0 1 2621
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1666464484
transform 1 0 2701 0 1 4665
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1666464484
transform 1 0 3151 0 1 4722
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1666464484
transform 1 0 2287 0 1 4722
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1666464484
transform 1 0 3050 0 1 6225
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1666464484
transform 1 0 3623 0 1 4722
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1666464484
transform 1 0 3722 0 1 6225
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1666464484
transform 1 0 4040 0 1 4665
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1666464484
transform 1 0 4418 0 1 4722
box 0 -1 93 308
use via1_2_x2_R90_512x8m81  via1_2_x2_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 3259 1 0 7937
box 0 -1 93 308
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_0
timestamp 1666464484
transform 0 1 4262 -1 0 544
box -1 -1 96 308
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_1
timestamp 1666464484
transform 0 1 2723 -1 0 544
box -1 -1 96 308
use via1_2_x2_R270_512x8m81  via1_2_x2_R270_512x8m81_2
timestamp 1666464484
transform 0 1 3182 -1 0 544
box -1 -1 96 308
use via1_512x8m81  via1_512x8m81_0
timestamp 1666464484
transform 1 0 3388 0 -1 6790
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 4506 1 0 3149
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_1
timestamp 1666464484
transform 0 -1 2486 1 0 3149
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_2
timestamp 1666464484
transform 0 -1 2520 1 0 4226
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_3
timestamp 1666464484
transform 0 -1 4396 1 0 4437
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_4
timestamp 1666464484
transform 0 -1 4568 1 0 4226
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_5
timestamp 1666464484
transform 0 -1 3595 1 0 5792
box 0 0 1 1
use via1_R90_512x8m81  via1_R90_512x8m81_6
timestamp 1666464484
transform 0 1 3276 1 0 5964
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_0
timestamp 1666464484
transform 0 -1 2925 -1 0 6762
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_1
timestamp 1666464484
transform 0 1 3083 -1 0 4321
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_2
timestamp 1666464484
transform 0 1 3193 -1 0 4532
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_3
timestamp 1666464484
transform 0 -1 3500 -1 0 7361
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_4
timestamp 1666464484
transform 0 -1 4060 -1 0 6740
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_5
timestamp 1666464484
transform 0 1 3659 -1 0 4321
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_6
timestamp 1666464484
transform 0 1 3371 -1 0 4321
box 0 0 1 1
use via1_R270_512x8m81  via1_R270_512x8m81_7
timestamp 1666464484
transform 0 1 3549 -1 0 4532
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1666464484
transform -1 0 4153 0 1 1018
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_1
timestamp 1666464484
transform 1 0 4276 0 1 1712
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_2
timestamp 1666464484
transform 1 0 3601 0 1 1018
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_3
timestamp 1666464484
transform -1 0 3920 0 1 1712
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_4
timestamp 1666464484
transform -1 0 3478 0 1 1712
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_5
timestamp 1666464484
transform 1 0 2596 0 1 6146
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_6
timestamp 1666464484
transform 1 0 4181 0 1 6146
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_7
timestamp 1666464484
transform 1 0 3503 0 1 6146
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_8
timestamp 1666464484
transform -1 0 3369 0 1 6146
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 4559 1 0 1494
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_1
timestamp 1666464484
transform 0 -1 3057 1 0 1505
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_2
timestamp 1666464484
transform 0 -1 3015 1 0 7728
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_3
timestamp 1666464484
transform 0 -1 2633 1 0 7937
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_4
timestamp 1666464484
transform 0 -1 3819 1 0 7728
box 0 0 1 1
use via1_x2_R90_512x8m81  via1_x2_R90_512x8m81_5
timestamp 1666464484
transform 0 -1 4497 1 0 7937
box 0 0 1 1
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_0
timestamp 1666464484
transform 0 1 2684 -1 0 4532
box 0 0 1 1
use via1_x2_R270_512x8m81  via1_x2_R270_512x8m81_1
timestamp 1666464484
transform 0 1 3883 -1 0 4532
box 0 0 1 1
use via2_x2_R90_512x8m81  via2_x2_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 1992 1 0 7728
box 0 0 1 1
<< labels >>
rlabel metal3 s 1179 5153 1179 5153 4 vdd
port 1 nsew
rlabel metal3 s 1247 2410 1247 2410 4 vss
port 2 nsew
rlabel metal3 s 1032 116 1032 116 4 vdd
port 1 nsew
rlabel metal2 s 3648 -136 3648 -136 4 qp
port 3 nsew
rlabel metal2 s 3995 7030 3995 7030 4 db
port 4 nsew
rlabel metal2 s 2868 7030 2868 7030 4 d
port 5 nsew
rlabel metal2 s 4111 -136 4111 -136 4 qn
port 6 nsew
rlabel metal1 s 3452 7551 3452 7551 4 wep
port 7 nsew
rlabel metal1 s 3437 7996 3437 7996 4 db
port 4 nsew
rlabel metal1 s 4471 2403 4471 2403 4 se
port 8 nsew
rlabel metal1 s 2040 7295 2040 7295 4 pcb
port 9 nsew
rlabel metal1 s 3432 7780 3432 7780 4 d
port 5 nsew
<< properties >>
string GDS_END 449718
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 435742
<< end >>
