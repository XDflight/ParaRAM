magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< ndiff >>
rect -1840 209 1840 228
rect -1840 163 -1821 209
rect -1775 163 -1697 209
rect -1651 163 -1573 209
rect -1527 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1527 209
rect 1573 163 1651 209
rect 1697 163 1775 209
rect 1821 163 1840 209
rect -1840 85 1840 163
rect -1840 39 -1821 85
rect -1775 39 -1697 85
rect -1651 39 -1573 85
rect -1527 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1527 85
rect 1573 39 1651 85
rect 1697 39 1775 85
rect 1821 39 1840 85
rect -1840 -39 1840 39
rect -1840 -85 -1821 -39
rect -1775 -85 -1697 -39
rect -1651 -85 -1573 -39
rect -1527 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1527 -39
rect 1573 -85 1651 -39
rect 1697 -85 1775 -39
rect 1821 -85 1840 -39
rect -1840 -163 1840 -85
rect -1840 -209 -1821 -163
rect -1775 -209 -1697 -163
rect -1651 -209 -1573 -163
rect -1527 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1527 -163
rect 1573 -209 1651 -163
rect 1697 -209 1775 -163
rect 1821 -209 1840 -163
rect -1840 -228 1840 -209
<< ndiffc >>
rect -1821 163 -1775 209
rect -1697 163 -1651 209
rect -1573 163 -1527 209
rect -1449 163 -1403 209
rect -1325 163 -1279 209
rect -1201 163 -1155 209
rect -1077 163 -1031 209
rect -953 163 -907 209
rect -829 163 -783 209
rect -705 163 -659 209
rect -581 163 -535 209
rect -457 163 -411 209
rect -333 163 -287 209
rect -209 163 -163 209
rect -85 163 -39 209
rect 39 163 85 209
rect 163 163 209 209
rect 287 163 333 209
rect 411 163 457 209
rect 535 163 581 209
rect 659 163 705 209
rect 783 163 829 209
rect 907 163 953 209
rect 1031 163 1077 209
rect 1155 163 1201 209
rect 1279 163 1325 209
rect 1403 163 1449 209
rect 1527 163 1573 209
rect 1651 163 1697 209
rect 1775 163 1821 209
rect -1821 39 -1775 85
rect -1697 39 -1651 85
rect -1573 39 -1527 85
rect -1449 39 -1403 85
rect -1325 39 -1279 85
rect -1201 39 -1155 85
rect -1077 39 -1031 85
rect -953 39 -907 85
rect -829 39 -783 85
rect -705 39 -659 85
rect -581 39 -535 85
rect -457 39 -411 85
rect -333 39 -287 85
rect -209 39 -163 85
rect -85 39 -39 85
rect 39 39 85 85
rect 163 39 209 85
rect 287 39 333 85
rect 411 39 457 85
rect 535 39 581 85
rect 659 39 705 85
rect 783 39 829 85
rect 907 39 953 85
rect 1031 39 1077 85
rect 1155 39 1201 85
rect 1279 39 1325 85
rect 1403 39 1449 85
rect 1527 39 1573 85
rect 1651 39 1697 85
rect 1775 39 1821 85
rect -1821 -85 -1775 -39
rect -1697 -85 -1651 -39
rect -1573 -85 -1527 -39
rect -1449 -85 -1403 -39
rect -1325 -85 -1279 -39
rect -1201 -85 -1155 -39
rect -1077 -85 -1031 -39
rect -953 -85 -907 -39
rect -829 -85 -783 -39
rect -705 -85 -659 -39
rect -581 -85 -535 -39
rect -457 -85 -411 -39
rect -333 -85 -287 -39
rect -209 -85 -163 -39
rect -85 -85 -39 -39
rect 39 -85 85 -39
rect 163 -85 209 -39
rect 287 -85 333 -39
rect 411 -85 457 -39
rect 535 -85 581 -39
rect 659 -85 705 -39
rect 783 -85 829 -39
rect 907 -85 953 -39
rect 1031 -85 1077 -39
rect 1155 -85 1201 -39
rect 1279 -85 1325 -39
rect 1403 -85 1449 -39
rect 1527 -85 1573 -39
rect 1651 -85 1697 -39
rect 1775 -85 1821 -39
rect -1821 -209 -1775 -163
rect -1697 -209 -1651 -163
rect -1573 -209 -1527 -163
rect -1449 -209 -1403 -163
rect -1325 -209 -1279 -163
rect -1201 -209 -1155 -163
rect -1077 -209 -1031 -163
rect -953 -209 -907 -163
rect -829 -209 -783 -163
rect -705 -209 -659 -163
rect -581 -209 -535 -163
rect -457 -209 -411 -163
rect -333 -209 -287 -163
rect -209 -209 -163 -163
rect -85 -209 -39 -163
rect 39 -209 85 -163
rect 163 -209 209 -163
rect 287 -209 333 -163
rect 411 -209 457 -163
rect 535 -209 581 -163
rect 659 -209 705 -163
rect 783 -209 829 -163
rect 907 -209 953 -163
rect 1031 -209 1077 -163
rect 1155 -209 1201 -163
rect 1279 -209 1325 -163
rect 1403 -209 1449 -163
rect 1527 -209 1573 -163
rect 1651 -209 1697 -163
rect 1775 -209 1821 -163
<< metal1 >>
rect -1832 209 1832 220
rect -1832 163 -1821 209
rect -1775 163 -1697 209
rect -1651 163 -1573 209
rect -1527 163 -1449 209
rect -1403 163 -1325 209
rect -1279 163 -1201 209
rect -1155 163 -1077 209
rect -1031 163 -953 209
rect -907 163 -829 209
rect -783 163 -705 209
rect -659 163 -581 209
rect -535 163 -457 209
rect -411 163 -333 209
rect -287 163 -209 209
rect -163 163 -85 209
rect -39 163 39 209
rect 85 163 163 209
rect 209 163 287 209
rect 333 163 411 209
rect 457 163 535 209
rect 581 163 659 209
rect 705 163 783 209
rect 829 163 907 209
rect 953 163 1031 209
rect 1077 163 1155 209
rect 1201 163 1279 209
rect 1325 163 1403 209
rect 1449 163 1527 209
rect 1573 163 1651 209
rect 1697 163 1775 209
rect 1821 163 1832 209
rect -1832 85 1832 163
rect -1832 39 -1821 85
rect -1775 39 -1697 85
rect -1651 39 -1573 85
rect -1527 39 -1449 85
rect -1403 39 -1325 85
rect -1279 39 -1201 85
rect -1155 39 -1077 85
rect -1031 39 -953 85
rect -907 39 -829 85
rect -783 39 -705 85
rect -659 39 -581 85
rect -535 39 -457 85
rect -411 39 -333 85
rect -287 39 -209 85
rect -163 39 -85 85
rect -39 39 39 85
rect 85 39 163 85
rect 209 39 287 85
rect 333 39 411 85
rect 457 39 535 85
rect 581 39 659 85
rect 705 39 783 85
rect 829 39 907 85
rect 953 39 1031 85
rect 1077 39 1155 85
rect 1201 39 1279 85
rect 1325 39 1403 85
rect 1449 39 1527 85
rect 1573 39 1651 85
rect 1697 39 1775 85
rect 1821 39 1832 85
rect -1832 -39 1832 39
rect -1832 -85 -1821 -39
rect -1775 -85 -1697 -39
rect -1651 -85 -1573 -39
rect -1527 -85 -1449 -39
rect -1403 -85 -1325 -39
rect -1279 -85 -1201 -39
rect -1155 -85 -1077 -39
rect -1031 -85 -953 -39
rect -907 -85 -829 -39
rect -783 -85 -705 -39
rect -659 -85 -581 -39
rect -535 -85 -457 -39
rect -411 -85 -333 -39
rect -287 -85 -209 -39
rect -163 -85 -85 -39
rect -39 -85 39 -39
rect 85 -85 163 -39
rect 209 -85 287 -39
rect 333 -85 411 -39
rect 457 -85 535 -39
rect 581 -85 659 -39
rect 705 -85 783 -39
rect 829 -85 907 -39
rect 953 -85 1031 -39
rect 1077 -85 1155 -39
rect 1201 -85 1279 -39
rect 1325 -85 1403 -39
rect 1449 -85 1527 -39
rect 1573 -85 1651 -39
rect 1697 -85 1775 -39
rect 1821 -85 1832 -39
rect -1832 -163 1832 -85
rect -1832 -209 -1821 -163
rect -1775 -209 -1697 -163
rect -1651 -209 -1573 -163
rect -1527 -209 -1449 -163
rect -1403 -209 -1325 -163
rect -1279 -209 -1201 -163
rect -1155 -209 -1077 -163
rect -1031 -209 -953 -163
rect -907 -209 -829 -163
rect -783 -209 -705 -163
rect -659 -209 -581 -163
rect -535 -209 -457 -163
rect -411 -209 -333 -163
rect -287 -209 -209 -163
rect -163 -209 -85 -163
rect -39 -209 39 -163
rect 85 -209 163 -163
rect 209 -209 287 -163
rect 333 -209 411 -163
rect 457 -209 535 -163
rect 581 -209 659 -163
rect 705 -209 783 -163
rect 829 -209 907 -163
rect 953 -209 1031 -163
rect 1077 -209 1155 -163
rect 1201 -209 1279 -163
rect 1325 -209 1403 -163
rect 1449 -209 1527 -163
rect 1573 -209 1651 -163
rect 1697 -209 1775 -163
rect 1821 -209 1832 -163
rect -1832 -220 1832 -209
<< properties >>
string GDS_END 830170
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 822294
<< end >>
