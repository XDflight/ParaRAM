magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 2464 844
rect 297 657 365 724
rect 1313 635 1537 724
rect 1471 506 1537 635
rect 1684 468 1730 676
rect 1888 514 1934 724
rect 2122 468 2236 676
rect 2326 506 2372 724
rect 1684 421 2236 468
rect 186 240 672 320
rect 2122 243 2236 421
rect 1674 192 2236 243
rect 317 60 385 127
rect 1344 60 1390 138
rect 1674 106 1720 192
rect 1887 60 1955 127
rect 2122 110 2236 192
rect 2346 60 2392 223
rect 0 -60 2464 60
<< obsm1 >>
rect 49 481 117 621
rect 49 413 653 481
rect 49 180 95 413
rect 744 382 790 632
rect 908 493 954 632
rect 908 447 1231 493
rect 744 336 1097 382
rect 1167 371 1231 447
rect 49 134 117 180
rect 744 154 821 336
rect 1167 325 2072 371
rect 1167 211 1231 325
rect 908 143 1231 211
<< labels >>
rlabel metal1 s 186 240 672 320 6 I
port 1 nsew default input
rlabel metal1 s 2122 468 2236 676 6 Z
port 2 nsew default output
rlabel metal1 s 1684 468 1730 676 6 Z
port 2 nsew default output
rlabel metal1 s 1684 421 2236 468 6 Z
port 2 nsew default output
rlabel metal1 s 2122 243 2236 421 6 Z
port 2 nsew default output
rlabel metal1 s 1674 192 2236 243 6 Z
port 2 nsew default output
rlabel metal1 s 2122 110 2236 192 6 Z
port 2 nsew default output
rlabel metal1 s 1674 110 1720 192 6 Z
port 2 nsew default output
rlabel metal1 s 1674 106 1720 110 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 2464 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 657 2372 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 657 1934 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 657 1537 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 635 2372 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 635 1934 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1313 635 1537 657 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 514 2372 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1888 514 1934 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1471 514 1537 635 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2326 506 2372 514 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1471 506 1537 514 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2346 138 2392 223 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2346 127 2392 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1344 127 1390 138 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2346 60 2392 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1887 60 1955 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1344 60 1390 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1083364
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1078096
<< end >>
