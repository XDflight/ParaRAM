magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 192
<< mvndiff >>
rect -88 179 0 192
rect -88 133 -75 179
rect -29 133 0 179
rect -88 59 0 133
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 179 208 192
rect 120 133 149 179
rect 195 133 208 179
rect 120 59 208 133
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 133 -29 179
rect -75 13 -29 59
rect 149 133 195 179
rect 149 13 195 59
<< polysilicon >>
rect 0 192 120 236
rect 0 -44 120 0
<< metal1 >>
rect -75 179 -29 192
rect -75 59 -29 133
rect -75 0 -29 13
rect 149 179 195 192
rect 149 59 195 133
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 96 -52 96 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 96 172 96 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 48704
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 47552
<< end >>
