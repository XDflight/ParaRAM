magic
tech gf180mcuC
timestamp 1666464484
<< properties >>
string GDS_END 2529370
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2529110
<< end >>
