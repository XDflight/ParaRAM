magic
tech gf180mcuC
timestamp 1666464484
<< metal1 >>
rect 0 111 316 123
rect 28 70 33 111
rect 45 65 50 104
rect 62 70 67 111
rect 79 65 84 104
rect 96 70 101 111
rect 113 65 118 104
rect 130 70 135 111
rect 147 65 152 104
rect 164 70 169 111
rect 181 65 186 104
rect 198 70 203 111
rect 215 65 220 104
rect 232 70 237 111
rect 249 65 254 104
rect 266 70 271 111
rect 283 76 288 104
rect 281 70 291 76
rect 300 70 305 111
rect 283 65 288 70
rect 45 59 288 65
rect 21 44 31 50
rect 45 47 50 59
rect 79 47 84 59
rect 113 47 118 59
rect 147 47 152 59
rect 181 47 186 59
rect 215 47 220 59
rect 249 47 254 59
rect 283 47 288 59
rect 45 41 288 47
rect 28 12 33 36
rect 45 19 50 41
rect 62 12 67 36
rect 79 19 84 41
rect 96 12 101 36
rect 113 19 118 41
rect 130 12 135 36
rect 147 19 152 41
rect 164 12 169 36
rect 181 19 186 41
rect 198 12 203 36
rect 215 19 220 41
rect 232 12 237 36
rect 249 19 254 41
rect 266 12 271 36
rect 283 19 288 41
rect 300 12 305 36
rect 0 0 316 12
<< obsm1 >>
rect 11 65 16 104
rect 11 59 40 65
rect 11 19 16 59
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 178 118 186 119
rect 202 118 210 119
rect 226 118 234 119
rect 250 118 258 119
rect 274 118 282 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 177 112 187 118
rect 201 112 211 118
rect 225 112 235 118
rect 249 112 259 118
rect 273 112 283 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 178 111 186 112
rect 202 111 210 112
rect 226 111 234 112
rect 250 111 258 112
rect 274 111 282 112
rect 281 69 291 77
rect 22 50 30 51
rect 21 44 31 50
rect 22 43 30 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 274 11 282 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 273 5 283 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
rect 274 4 282 5
<< labels >>
rlabel metal2 s 22 43 30 51 6 A
port 1 nsew signal input
rlabel metal2 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal1 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 178 111 186 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 177 112 187 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 202 111 210 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 201 112 211 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 226 111 234 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 225 112 235 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 250 111 258 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 249 112 259 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 274 111 282 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 273 112 283 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 28 70 33 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 62 70 67 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 96 70 101 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 130 70 135 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 164 70 169 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 198 70 203 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 232 70 237 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 266 70 271 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 300 70 305 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 111 316 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 274 4 282 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 273 5 283 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 62 0 67 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 96 0 101 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 130 0 135 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 164 0 169 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 198 0 203 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 232 0 237 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 266 0 271 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 300 0 305 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 316 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 281 69 291 77 6 Y
port 4 nsew signal output
rlabel metal1 s 45 19 50 104 6 Y
port 4 nsew signal output
rlabel metal1 s 79 19 84 104 6 Y
port 4 nsew signal output
rlabel metal1 s 113 19 118 104 6 Y
port 4 nsew signal output
rlabel metal1 s 147 19 152 104 6 Y
port 4 nsew signal output
rlabel metal1 s 181 19 186 104 6 Y
port 4 nsew signal output
rlabel metal1 s 215 19 220 104 6 Y
port 4 nsew signal output
rlabel metal1 s 249 19 254 104 6 Y
port 4 nsew signal output
rlabel metal1 s 45 41 288 47 6 Y
port 4 nsew signal output
rlabel metal1 s 45 59 288 65 6 Y
port 4 nsew signal output
rlabel metal1 s 283 19 288 104 6 Y
port 4 nsew signal output
rlabel metal1 s 281 70 291 76 6 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 316 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
