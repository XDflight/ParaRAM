magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 322
<< polysilicon >>
rect -31 191 88 222
rect -30 -73 88 0
use pmos_5p04310591302041_512x8m81  pmos_5p04310591302041_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 312
<< properties >>
string GDS_END 61726
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 61412
<< end >>
