magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 522 88 595
rect 193 522 312 595
rect -31 -74 88 -1
rect 193 -74 312 -1
use nmos_5p04310591302029_512x8m81  nmos_5p04310591302029_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 432 566
<< properties >>
string GDS_END 336070
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 335692
<< end >>
