magic
tech gf180mcuC
timestamp 1666464484
<< metal1 >>
rect -155 150 25 162
rect -126 125 -121 150
rect -58 109 -53 150
rect -118 83 -108 89
rect -86 83 -76 89
rect -51 83 -41 89
rect -9 109 -4 150
rect 8 103 13 143
rect 8 102 16 103
rect -126 12 -118 36
rect 8 96 18 102
rect 8 95 16 96
rect -61 12 -53 36
rect -9 12 -4 36
rect 8 19 13 95
rect -155 0 25 12
<< obsm1 >>
rect -143 77 -138 143
rect -92 114 -87 143
rect -132 109 -87 114
rect -41 110 -36 143
rect -132 89 -127 109
rect -41 105 -31 110
rect -103 94 -93 100
rect -133 83 -124 89
rect -145 76 -138 77
rect -148 70 -138 76
rect -146 69 -138 70
rect -143 19 -138 69
rect -132 46 -127 83
rect -101 57 -95 94
rect -65 70 -55 76
rect -36 57 -31 105
rect -26 106 -21 143
rect -26 102 -18 106
rect -26 101 -16 102
rect -26 96 1 101
rect -26 95 -18 96
rect -20 70 -10 76
rect -101 51 -31 57
rect -132 41 -87 46
rect -36 44 -31 51
rect -5 46 1 96
rect -92 19 -87 41
rect -41 39 -31 44
rect -26 41 1 46
rect -41 19 -36 39
rect -26 19 -21 41
<< metal2 >>
rect -145 157 -137 158
rect -121 157 -113 158
rect -97 157 -89 158
rect -73 157 -65 158
rect -49 157 -41 158
rect -25 157 -17 158
rect -1 157 7 158
rect -146 151 -136 157
rect -122 151 -112 157
rect -98 151 -88 157
rect -74 151 -64 157
rect -50 151 -40 157
rect -26 151 -16 157
rect -2 151 8 157
rect -145 150 -137 151
rect -121 150 -113 151
rect -97 150 -89 151
rect -73 150 -65 151
rect -49 150 -41 151
rect -25 150 -17 151
rect -1 150 7 151
rect 9 102 17 103
rect 8 96 18 102
rect 9 95 17 96
rect -118 82 -108 90
rect -85 89 -77 90
rect -51 89 -41 90
rect -86 83 -41 89
rect -85 82 -77 83
rect -51 82 -41 83
rect -145 11 -137 12
rect -121 11 -113 12
rect -97 11 -89 12
rect -73 11 -65 12
rect -49 11 -41 12
rect -25 11 -17 12
rect -1 11 7 12
rect -146 5 -136 11
rect -122 5 -112 11
rect -98 5 -88 11
rect -74 5 -64 11
rect -50 5 -40 11
rect -26 5 -16 11
rect -2 5 8 11
rect -145 4 -137 5
rect -121 4 -113 5
rect -97 4 -89 5
rect -73 4 -65 5
rect -49 4 -41 5
rect -25 4 -17 5
rect -1 4 7 5
<< obsm2 >>
rect -25 102 -17 103
rect -26 96 -16 102
rect -25 95 -17 96
rect -148 76 -138 77
rect -64 76 -56 77
rect -20 76 -10 77
rect -148 70 -10 76
rect -148 69 -138 70
rect -64 69 -56 70
rect -20 69 -10 70
<< labels >>
rlabel metal2 s -85 82 -77 90 4 CLKN
port 1 nsew clock input
rlabel metal2 s -86 83 -41 89 4 CLKN
port 1 nsew clock input
rlabel metal2 s -51 82 -41 90 4 CLKN
port 1 nsew clock input
rlabel metal1 s -86 83 -76 89 4 CLKN
port 1 nsew clock input
rlabel metal1 s -51 83 -41 89 4 CLKN
port 1 nsew clock input
rlabel metal2 s -118 82 -108 90 4 D
port 2 nsew signal input
rlabel metal1 s -118 83 -108 89 4 D
port 2 nsew signal input
rlabel metal2 s 9 95 17 103 6 Q
port 3 nsew signal output
rlabel metal2 s 8 96 18 102 6 Q
port 3 nsew signal output
rlabel metal1 s 8 19 13 143 6 Q
port 3 nsew signal output
rlabel metal1 s 8 95 16 103 6 Q
port 3 nsew signal output
rlabel metal1 s 8 96 18 102 6 Q
port 3 nsew signal output
rlabel metal2 s -145 150 -137 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -146 151 -136 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -121 150 -113 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -122 151 -112 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -97 150 -89 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -98 151 -88 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -73 150 -65 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -74 151 -64 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -49 150 -41 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -50 151 -40 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -25 150 -17 158 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -26 151 -16 157 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -1 150 7 158 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -2 151 8 157 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s -126 125 -121 162 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s -58 109 -53 162 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s -9 109 -4 162 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s -155 150 25 162 4 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s -145 4 -137 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -146 5 -136 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -121 4 -113 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -122 5 -112 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -97 4 -89 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -98 5 -88 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -73 4 -65 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -74 5 -64 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -49 4 -41 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -50 5 -40 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -25 4 -17 12 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -26 5 -16 11 4 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -1 4 7 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s -2 5 8 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s -126 0 -118 36 4 VSS
port 5 nsew ground bidirectional
rlabel metal1 s -61 0 -53 36 4 VSS
port 5 nsew ground bidirectional
rlabel metal1 s -9 0 -4 36 4 VSS
port 5 nsew ground bidirectional
rlabel metal1 s -155 0 25 12 4 VSS
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX -155 0 25 162
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
