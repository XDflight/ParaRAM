magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 1344 844
rect 132 217 204 574
rect 356 316 452 656
rect 580 316 676 656
rect 804 316 900 656
rect 1017 506 1063 724
rect 38 60 106 152
rect 522 60 590 152
rect 1017 60 1063 171
rect 1214 126 1315 676
rect 0 -60 1344 60
<< obsm1 >>
rect 56 624 306 670
rect 260 266 306 624
rect 1103 266 1153 454
rect 260 219 1153 266
rect 298 106 366 219
rect 746 106 814 219
<< labels >>
rlabel metal1 s 132 217 204 574 6 A1
port 1 nsew default input
rlabel metal1 s 356 316 452 656 6 A2
port 2 nsew default input
rlabel metal1 s 580 316 676 656 6 A3
port 3 nsew default input
rlabel metal1 s 804 316 900 656 6 A4
port 4 nsew default input
rlabel metal1 s 1214 126 1315 676 6 Z
port 5 nsew default output
rlabel metal1 s 0 724 1344 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1017 506 1063 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1017 152 1063 171 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1017 60 1063 152 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 522 60 590 152 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 152 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1344 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 167626
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 163996
<< end >>
