magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 1362
<< mvndiff >>
rect -88 1349 0 1362
rect -88 1303 -75 1349
rect -29 1303 0 1349
rect -88 1242 0 1303
rect -88 1196 -75 1242
rect -29 1196 0 1242
rect -88 1135 0 1196
rect -88 1089 -75 1135
rect -29 1089 0 1135
rect -88 1028 0 1089
rect -88 982 -75 1028
rect -29 982 0 1028
rect -88 921 0 982
rect -88 875 -75 921
rect -29 875 0 921
rect -88 814 0 875
rect -88 768 -75 814
rect -29 768 0 814
rect -88 707 0 768
rect -88 661 -75 707
rect -29 661 0 707
rect -88 599 0 661
rect -88 553 -75 599
rect -29 553 0 599
rect -88 491 0 553
rect -88 445 -75 491
rect -29 445 0 491
rect -88 383 0 445
rect -88 337 -75 383
rect -29 337 0 383
rect -88 275 0 337
rect -88 229 -75 275
rect -29 229 0 275
rect -88 167 0 229
rect -88 121 -75 167
rect -29 121 0 167
rect -88 59 0 121
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1349 208 1362
rect 120 1303 149 1349
rect 195 1303 208 1349
rect 120 1242 208 1303
rect 120 1196 149 1242
rect 195 1196 208 1242
rect 120 1135 208 1196
rect 120 1089 149 1135
rect 195 1089 208 1135
rect 120 1028 208 1089
rect 120 982 149 1028
rect 195 982 208 1028
rect 120 921 208 982
rect 120 875 149 921
rect 195 875 208 921
rect 120 814 208 875
rect 120 768 149 814
rect 195 768 208 814
rect 120 707 208 768
rect 120 661 149 707
rect 195 661 208 707
rect 120 599 208 661
rect 120 553 149 599
rect 195 553 208 599
rect 120 491 208 553
rect 120 445 149 491
rect 195 445 208 491
rect 120 383 208 445
rect 120 337 149 383
rect 195 337 208 383
rect 120 275 208 337
rect 120 229 149 275
rect 195 229 208 275
rect 120 167 208 229
rect 120 121 149 167
rect 195 121 208 167
rect 120 59 208 121
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 1303 -29 1349
rect -75 1196 -29 1242
rect -75 1089 -29 1135
rect -75 982 -29 1028
rect -75 875 -29 921
rect -75 768 -29 814
rect -75 661 -29 707
rect -75 553 -29 599
rect -75 445 -29 491
rect -75 337 -29 383
rect -75 229 -29 275
rect -75 121 -29 167
rect -75 13 -29 59
rect 149 1303 195 1349
rect 149 1196 195 1242
rect 149 1089 195 1135
rect 149 982 195 1028
rect 149 875 195 921
rect 149 768 195 814
rect 149 661 195 707
rect 149 553 195 599
rect 149 445 195 491
rect 149 337 195 383
rect 149 229 195 275
rect 149 121 195 167
rect 149 13 195 59
<< polysilicon >>
rect 0 1362 120 1406
rect 0 -44 120 0
<< metal1 >>
rect -75 1349 -29 1362
rect -75 1242 -29 1303
rect -75 1135 -29 1196
rect -75 1028 -29 1089
rect -75 921 -29 982
rect -75 814 -29 875
rect -75 707 -29 768
rect -75 599 -29 661
rect -75 491 -29 553
rect -75 383 -29 445
rect -75 275 -29 337
rect -75 167 -29 229
rect -75 59 -29 121
rect -75 0 -29 13
rect 149 1349 195 1362
rect 149 1242 195 1303
rect 149 1135 195 1196
rect 149 1028 195 1089
rect 149 921 195 982
rect 149 814 195 875
rect 149 707 195 768
rect 149 599 195 661
rect 149 491 195 553
rect 149 383 195 445
rect 149 275 195 337
rect 149 167 195 229
rect 149 59 195 121
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 681 -52 681 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 681 172 681 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 15252
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 12692
<< end >>
