magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 4071 10025 5372 10041
rect 3785 9887 5372 10025
rect 3785 9377 6659 9887
rect 3785 9364 5372 9377
rect 3787 7478 4285 7496
rect 3582 3757 4285 7478
rect 5326 4684 5539 7477
rect 4812 4661 5539 4684
rect 5967 4662 7077 7575
rect 5432 1986 5434 1987
rect 5432 797 5500 1986
<< pmos >>
rect 4326 9505 4446 9846
rect 4549 9505 4669 9846
rect 4774 9505 4894 9846
rect 4997 9505 5117 9846
<< pdiff >>
rect 4207 9801 4326 9846
rect 4207 9755 4251 9801
rect 4297 9755 4326 9801
rect 4207 9597 4326 9755
rect 4207 9551 4251 9597
rect 4297 9551 4326 9597
rect 4207 9505 4326 9551
rect 4446 9505 4549 9846
rect 4669 9801 4774 9846
rect 4669 9755 4699 9801
rect 4745 9755 4774 9801
rect 4669 9597 4774 9755
rect 4669 9551 4699 9597
rect 4745 9551 4774 9597
rect 4669 9505 4774 9551
rect 4894 9505 4997 9846
rect 5117 9801 5236 9846
rect 5117 9755 5147 9801
rect 5193 9755 5236 9801
rect 5117 9597 5236 9755
rect 5117 9551 5147 9597
rect 5193 9551 5236 9597
rect 5117 9505 5236 9551
<< pdiffc >>
rect 4251 9755 4297 9801
rect 4251 9551 4297 9597
rect 4699 9755 4745 9801
rect 4699 9551 4745 9597
rect 5147 9755 5193 9801
rect 5147 9551 5193 9597
<< nsubdiff >>
rect 3948 9797 4032 9816
rect 3948 9563 3967 9797
rect 4013 9563 4032 9797
rect 3948 9544 4032 9563
rect 6440 9797 6524 9816
rect 6440 9563 6459 9797
rect 6505 9563 6524 9797
rect 6440 9544 6524 9563
rect 3728 7170 4011 7330
<< nsubdiffcont >>
rect 3967 9563 4013 9797
rect 6459 9563 6505 9797
<< polysilicon >>
rect 4550 10512 4669 10513
rect 4886 10445 4970 10464
rect 4886 10305 4905 10445
rect 4951 10305 4970 10445
rect 4550 10209 4669 10239
rect 4326 10121 4446 10209
rect 4550 10180 4670 10209
rect 4886 10180 4970 10305
rect 4550 10167 4970 10180
rect 4153 10102 4446 10121
rect 4153 10056 4172 10102
rect 4312 10056 4446 10102
rect 4153 10037 4446 10056
rect 4326 9846 4446 10037
rect 4549 10074 4970 10167
rect 4549 9846 4669 10074
rect 4774 10063 4970 10074
rect 4774 9846 4894 10063
rect 5081 9993 5275 10051
rect 5081 9967 5100 9993
rect 4997 9947 5100 9967
rect 5240 9947 5275 9993
rect 4997 9907 5275 9947
rect 4997 9846 5117 9907
rect 5920 9882 6040 10205
rect 5802 9807 6146 9882
rect 5802 9746 5922 9807
rect 6026 9746 6146 9807
rect 4326 9432 4446 9505
rect 4549 9432 4669 9505
rect 4774 9432 4894 9505
rect 4997 9432 5117 9505
rect 5802 9459 5922 9497
rect 6026 9459 6146 9497
rect 5802 9440 6146 9459
rect 5802 9394 5868 9440
rect 6102 9394 6146 9440
rect 5802 9375 6146 9394
rect 173 3782 366 3827
rect 173 3736 247 3782
rect 293 3736 366 3782
rect 173 3690 366 3736
rect 1425 3782 1618 3827
rect 1425 3736 1499 3782
rect 1545 3736 1618 3782
rect 1425 3690 1618 3736
rect 1965 3578 2158 3623
rect 1965 3532 2039 3578
rect 2085 3532 2158 3578
rect 1965 3486 2158 3532
rect 3217 3578 3410 3623
rect 3217 3532 3291 3578
rect 3337 3532 3410 3578
rect 3217 3486 3410 3532
rect 397 3374 590 3419
rect 397 3328 471 3374
rect 517 3328 590 3374
rect 397 3282 590 3328
rect 2189 3374 2382 3419
rect 2189 3328 2263 3374
rect 2309 3328 2382 3374
rect 2189 3282 2382 3328
rect 1201 3174 1394 3219
rect 1201 3128 1275 3174
rect 1321 3128 1394 3174
rect 1201 3082 1394 3128
rect 2993 3174 3186 3219
rect 2993 3128 3067 3174
rect 3113 3128 3186 3174
rect 2993 3082 3186 3128
<< polycontact >>
rect 4905 10305 4951 10445
rect 4172 10056 4312 10102
rect 5100 9947 5240 9993
rect 5868 9394 6102 9440
rect 247 3736 293 3782
rect 1499 3736 1545 3782
rect 2039 3532 2085 3578
rect 3291 3532 3337 3578
rect 471 3328 517 3374
rect 2263 3328 2309 3374
rect 1275 3128 1321 3174
rect 3067 3128 3113 3174
<< metal1 >>
rect 4215 11315 4332 11393
rect 4215 10859 4331 11315
rect 4663 10859 4779 11399
rect 4203 10820 4331 10859
rect 4203 10768 4241 10820
rect 4293 10768 4331 10820
rect 4203 10602 4331 10768
rect 4203 10550 4241 10602
rect 4293 10550 4331 10602
rect 4642 10820 4779 10859
rect 4642 10768 4680 10820
rect 4732 10768 4779 10820
rect 6034 11315 6150 11433
rect 6034 10803 6149 11315
rect 6034 10802 6150 10803
rect 4642 10602 4779 10768
rect 6026 10763 6154 10802
rect 6026 10711 6064 10763
rect 6116 10711 6154 10763
rect 4203 10384 4331 10550
rect 4203 10332 4241 10384
rect 4293 10332 4331 10384
rect 4203 10292 4331 10332
rect 4215 10240 4331 10292
rect 4439 10152 4555 10554
rect 4642 10550 4680 10602
rect 4732 10550 4779 10602
rect 4642 10384 4779 10550
rect 4642 10332 4680 10384
rect 4732 10332 4779 10384
rect 4642 10292 4779 10332
rect 4864 10604 4988 10644
rect 4864 10552 4900 10604
rect 4952 10552 4988 10604
rect 4864 10445 4988 10552
rect 4864 10386 4905 10445
rect 4951 10386 4988 10445
rect 6026 10545 6154 10711
rect 6026 10493 6064 10545
rect 6116 10493 6154 10545
rect 4864 10334 4900 10386
rect 4952 10334 4988 10386
rect 4864 10305 4905 10334
rect 4951 10305 4988 10334
rect 4864 10294 4988 10305
rect 4663 10240 4779 10292
rect 4143 10102 4323 10114
rect 4143 10050 4155 10102
rect 4312 10056 4323 10102
rect 4311 10050 4323 10056
rect 4143 10038 4323 10050
rect 4439 10033 4779 10152
rect 5845 10121 5891 10417
rect 6026 10327 6154 10493
rect 6026 10275 6064 10327
rect 6116 10275 6154 10327
rect 6026 10235 6154 10275
rect 7060 10121 7184 10154
rect 5845 10114 7186 10121
rect 5071 10102 5251 10114
rect 5071 10050 5083 10102
rect 5239 10050 5251 10102
rect 5071 10038 5251 10050
rect 4215 9837 4331 9851
rect 3929 9797 4053 9837
rect 3929 9745 3965 9797
rect 4017 9745 4053 9797
rect 3929 9579 3967 9745
rect 4013 9579 4053 9745
rect 3929 9527 3965 9579
rect 4017 9527 4053 9579
rect 3929 9487 4053 9527
rect 4205 9801 4331 9837
rect 4205 9797 4251 9801
rect 4205 9745 4241 9797
rect 4297 9755 4331 9801
rect 4293 9745 4331 9755
rect 4205 9597 4331 9745
rect 4205 9579 4251 9597
rect 4205 9527 4241 9579
rect 4297 9551 4331 9597
rect 4293 9527 4331 9551
rect 4205 9514 4331 9527
rect 4663 9801 4779 10033
rect 5089 9993 5251 10038
rect 5089 9947 5100 9993
rect 5240 9947 5251 9993
rect 5845 10062 7096 10114
rect 7148 10062 7186 10114
rect 5845 9987 7186 10062
rect 5089 9936 5251 9947
rect 4663 9755 4699 9801
rect 4745 9755 4779 9801
rect 4663 9597 4779 9755
rect 4663 9551 4699 9597
rect 4745 9551 4779 9597
rect 4205 9487 4329 9514
rect 4663 9434 4779 9551
rect 5111 9801 5773 9851
rect 5111 9755 5147 9801
rect 5193 9755 5773 9801
rect 5111 9629 5773 9755
rect 5111 9597 5325 9629
rect 5111 9551 5147 9597
rect 5193 9577 5325 9597
rect 5377 9577 5537 9629
rect 5589 9577 5773 9629
rect 5951 9616 5997 9987
rect 7060 9896 7184 9987
rect 6175 9811 6545 9851
rect 6175 9759 6454 9811
rect 6506 9759 6545 9811
rect 7060 9844 7096 9896
rect 7148 9844 7184 9896
rect 7060 9804 7184 9844
rect 5193 9551 5773 9577
rect 5111 9519 5773 9551
rect 6175 9593 6459 9759
rect 6505 9593 6545 9759
rect 6175 9541 6454 9593
rect 6506 9541 6545 9593
rect 6175 9527 6545 9541
rect 5111 9514 5227 9519
rect 6418 9501 6542 9527
rect 5857 9440 6113 9451
rect 5857 9434 5868 9440
rect 4663 9394 5868 9434
rect 6102 9394 6113 9440
rect 4663 9393 6113 9394
rect 4663 9341 5323 9393
rect 5375 9341 5535 9393
rect 5587 9341 6113 9393
rect 4663 9314 6113 9341
rect 5285 9301 5625 9314
rect 4009 7309 4134 7310
rect 3627 7190 4134 7309
rect 212 3782 327 3818
rect 212 3736 247 3782
rect 293 3736 327 3782
rect 212 3699 327 3736
rect 1464 3782 1579 3818
rect 1464 3736 1499 3782
rect 1545 3736 1579 3782
rect 1464 3699 1579 3736
rect 4591 3710 4720 4256
rect 2004 3578 2119 3614
rect 2004 3532 2039 3578
rect 2085 3532 2119 3578
rect 2004 3495 2119 3532
rect 3256 3578 3371 3614
rect 3256 3532 3291 3578
rect 3337 3532 3371 3578
rect 3256 3495 3371 3532
rect 5105 3581 5234 3622
rect 5105 3529 5143 3581
rect 5195 3529 5234 3581
rect 5105 3488 5234 3529
rect 436 3374 551 3410
rect 436 3328 471 3374
rect 517 3328 551 3374
rect 436 3291 551 3328
rect 2228 3374 2343 3410
rect 2228 3328 2263 3374
rect 2309 3328 2343 3374
rect 2228 3291 2343 3328
rect 6282 3379 6411 3420
rect 6282 3327 6320 3379
rect 6372 3327 6411 3379
rect 6282 3286 6411 3327
rect 1240 3174 1355 3210
rect 1240 3128 1275 3174
rect 1321 3128 1355 3174
rect 1240 3091 1355 3128
rect 3032 3174 3147 3210
rect 3032 3128 3067 3174
rect 3113 3128 3147 3174
rect 3032 3091 3147 3128
rect 6796 3177 6925 3218
rect 6796 3125 6834 3177
rect 6886 3125 6925 3177
rect 6796 3084 6925 3125
<< via1 >>
rect 4241 10768 4293 10820
rect 4241 10550 4293 10602
rect 4680 10768 4732 10820
rect 6064 10711 6116 10763
rect 4241 10332 4293 10384
rect 4680 10550 4732 10602
rect 4680 10332 4732 10384
rect 4900 10552 4952 10604
rect 6064 10493 6116 10545
rect 4900 10334 4905 10386
rect 4905 10334 4951 10386
rect 4951 10334 4952 10386
rect 4155 10056 4172 10102
rect 4172 10056 4311 10102
rect 4155 10050 4311 10056
rect 6064 10275 6116 10327
rect 5083 10050 5239 10102
rect 3965 9745 3967 9797
rect 3967 9745 4013 9797
rect 4013 9745 4017 9797
rect 3965 9563 3967 9579
rect 3967 9563 4013 9579
rect 4013 9563 4017 9579
rect 3965 9527 4017 9563
rect 4241 9755 4251 9797
rect 4251 9755 4293 9797
rect 4241 9745 4293 9755
rect 4241 9551 4251 9579
rect 4251 9551 4293 9579
rect 4241 9527 4293 9551
rect 7096 10062 7148 10114
rect 5325 9577 5377 9629
rect 5537 9577 5589 9629
rect 6454 9797 6506 9811
rect 6454 9759 6459 9797
rect 6459 9759 6505 9797
rect 6505 9759 6506 9797
rect 7096 9844 7148 9896
rect 6454 9563 6459 9593
rect 6459 9563 6505 9593
rect 6505 9563 6506 9593
rect 6454 9541 6506 9563
rect 5323 9341 5375 9393
rect 5535 9341 5587 9393
rect 5143 3529 5195 3581
rect 6320 3327 6372 3379
rect 6834 3125 6886 3177
<< metal2 >>
rect 653 11057 783 11191
rect 1009 11057 1139 11191
rect 2443 11057 2573 11191
rect 2805 11057 2935 11191
rect 4203 10822 4331 10859
rect 4203 10766 4239 10822
rect 4295 10766 4331 10822
rect 4203 10604 4331 10766
rect 4203 10548 4239 10604
rect 4295 10548 4331 10604
rect 4203 10386 4331 10548
rect 4203 10330 4239 10386
rect 4295 10330 4331 10386
rect 4203 10292 4331 10330
rect 4642 10822 4770 10859
rect 4642 10766 4678 10822
rect 4734 10766 4770 10822
rect 4642 10604 4770 10766
rect 6026 10765 6154 10802
rect 6026 10709 6062 10765
rect 6118 10709 6154 10765
rect 4642 10548 4678 10604
rect 4734 10548 4770 10604
rect 4642 10386 4770 10548
rect 4861 10604 4990 10645
rect 4861 10552 4900 10604
rect 4952 10552 4990 10604
rect 4861 10511 4990 10552
rect 6026 10547 6154 10709
rect 4642 10330 4678 10386
rect 4734 10330 4770 10386
rect 4642 10292 4770 10330
rect 4864 10386 4988 10511
rect 4864 10334 4900 10386
rect 4952 10334 4988 10386
rect 4864 10294 4988 10334
rect 6026 10491 6062 10547
rect 6118 10491 6154 10547
rect 6026 10329 6154 10491
rect 6026 10273 6062 10329
rect 6118 10273 6154 10329
rect 6026 10235 6154 10273
rect 4013 10102 5251 10155
rect 4013 10050 4155 10102
rect 4311 10050 5083 10102
rect 5239 10050 5251 10102
rect 4013 10021 5251 10050
rect 7060 10114 7184 10154
rect 7060 10062 7096 10114
rect 7148 10062 7184 10114
rect 7060 9974 7184 10062
rect 7057 9896 7186 9974
rect 6418 9850 6542 9851
rect 3929 9836 4053 9837
rect 4205 9836 4329 9837
rect 3927 9799 4055 9836
rect 3927 9743 3963 9799
rect 4019 9743 4055 9799
rect 3927 9581 4055 9743
rect 3927 9525 3963 9581
rect 4019 9525 4055 9581
rect 3927 9363 4055 9525
rect 3927 9307 3963 9363
rect 4019 9307 4055 9363
rect 3927 9269 4055 9307
rect 4203 9799 4331 9836
rect 4203 9743 4239 9799
rect 4295 9743 4331 9799
rect 4203 9581 4331 9743
rect 6416 9813 6544 9850
rect 6416 9757 6452 9813
rect 6508 9757 6544 9813
rect 4203 9525 4239 9581
rect 4295 9525 4331 9581
rect 5287 9631 5627 9670
rect 5287 9575 5323 9631
rect 5379 9575 5535 9631
rect 5591 9575 5627 9631
rect 5287 9536 5627 9575
rect 6416 9595 6544 9757
rect 6416 9539 6452 9595
rect 6508 9539 6544 9595
rect 4203 9363 4331 9525
rect 4203 9307 4239 9363
rect 4295 9307 4331 9363
rect 4203 9269 4331 9307
rect 5286 9393 5625 9434
rect 5286 9341 5323 9393
rect 5375 9341 5535 9393
rect 5587 9341 5625 9393
rect 5286 9301 5625 9341
rect 6416 9377 6544 9539
rect 6416 9321 6452 9377
rect 6508 9321 6544 9377
rect 5390 9300 5520 9301
rect 5390 5473 5519 9300
rect 6416 9283 6544 9321
rect 7057 9844 7096 9896
rect 7148 9844 7186 9896
rect 4876 5340 5519 5473
rect 4876 3674 5005 5340
rect 5105 3581 5234 5163
rect 5105 3529 5143 3581
rect 5195 3529 5234 3581
rect 5105 3488 5234 3529
rect 6282 3379 6411 4256
rect 6282 3327 6320 3379
rect 6372 3327 6411 3379
rect 6282 3286 6411 3327
rect 6796 3177 6925 5163
rect 7057 4259 7186 9844
rect 6796 3125 6834 3177
rect 6886 3125 6925 3177
rect 6796 3084 6925 3125
rect 5160 212 5289 346
rect 6851 212 6980 346
<< via2 >>
rect 4239 10820 4295 10822
rect 4239 10768 4241 10820
rect 4241 10768 4293 10820
rect 4293 10768 4295 10820
rect 4239 10766 4295 10768
rect 4239 10602 4295 10604
rect 4239 10550 4241 10602
rect 4241 10550 4293 10602
rect 4293 10550 4295 10602
rect 4239 10548 4295 10550
rect 4239 10384 4295 10386
rect 4239 10332 4241 10384
rect 4241 10332 4293 10384
rect 4293 10332 4295 10384
rect 4239 10330 4295 10332
rect 4678 10820 4734 10822
rect 4678 10768 4680 10820
rect 4680 10768 4732 10820
rect 4732 10768 4734 10820
rect 4678 10766 4734 10768
rect 6062 10763 6118 10765
rect 6062 10711 6064 10763
rect 6064 10711 6116 10763
rect 6116 10711 6118 10763
rect 6062 10709 6118 10711
rect 4678 10602 4734 10604
rect 4678 10550 4680 10602
rect 4680 10550 4732 10602
rect 4732 10550 4734 10602
rect 4678 10548 4734 10550
rect 4678 10384 4734 10386
rect 4678 10332 4680 10384
rect 4680 10332 4732 10384
rect 4732 10332 4734 10384
rect 4678 10330 4734 10332
rect 6062 10545 6118 10547
rect 6062 10493 6064 10545
rect 6064 10493 6116 10545
rect 6116 10493 6118 10545
rect 6062 10491 6118 10493
rect 6062 10327 6118 10329
rect 6062 10275 6064 10327
rect 6064 10275 6116 10327
rect 6116 10275 6118 10327
rect 6062 10273 6118 10275
rect 3963 9797 4019 9799
rect 3963 9745 3965 9797
rect 3965 9745 4017 9797
rect 4017 9745 4019 9797
rect 3963 9743 4019 9745
rect 3963 9579 4019 9581
rect 3963 9527 3965 9579
rect 3965 9527 4017 9579
rect 4017 9527 4019 9579
rect 3963 9525 4019 9527
rect 3963 9307 4019 9363
rect 4239 9797 4295 9799
rect 4239 9745 4241 9797
rect 4241 9745 4293 9797
rect 4293 9745 4295 9797
rect 4239 9743 4295 9745
rect 6452 9811 6508 9813
rect 6452 9759 6454 9811
rect 6454 9759 6506 9811
rect 6506 9759 6508 9811
rect 6452 9757 6508 9759
rect 4239 9579 4295 9581
rect 4239 9527 4241 9579
rect 4241 9527 4293 9579
rect 4293 9527 4295 9579
rect 4239 9525 4295 9527
rect 5323 9629 5379 9631
rect 5323 9577 5325 9629
rect 5325 9577 5377 9629
rect 5377 9577 5379 9629
rect 5323 9575 5379 9577
rect 5535 9629 5591 9631
rect 5535 9577 5537 9629
rect 5537 9577 5589 9629
rect 5589 9577 5591 9629
rect 5535 9575 5591 9577
rect 6452 9593 6508 9595
rect 6452 9541 6454 9593
rect 6454 9541 6506 9593
rect 6506 9541 6508 9593
rect 6452 9539 6508 9541
rect 4239 9307 4295 9363
rect 6452 9321 6508 9377
<< metal3 >>
rect -289 10822 7380 10971
rect -289 10766 4239 10822
rect 4295 10766 4678 10822
rect 4734 10766 7380 10822
rect -289 10765 7380 10766
rect -289 10709 6062 10765
rect 6118 10709 7380 10765
rect -289 10604 7380 10709
rect -289 10548 4239 10604
rect 4295 10548 4678 10604
rect 4734 10548 7380 10604
rect -289 10547 7380 10548
rect -289 10491 6062 10547
rect 6118 10491 7380 10547
rect -289 10386 7380 10491
rect -289 10330 4239 10386
rect 4295 10330 4678 10386
rect 4734 10330 7380 10386
rect -289 10329 7380 10330
rect -289 10273 6062 10329
rect 6118 10273 7380 10329
rect -289 10019 7380 10273
rect -289 9813 7380 9907
rect -289 9799 6452 9813
rect -289 9743 3963 9799
rect 4019 9743 4239 9799
rect 4295 9757 6452 9799
rect 6508 9757 7380 9813
rect 4295 9743 7380 9757
rect -289 9631 7380 9743
rect -289 9581 5323 9631
rect -289 9525 3963 9581
rect 4019 9525 4239 9581
rect 4295 9575 5323 9581
rect 5379 9575 5535 9631
rect 5591 9595 7380 9631
rect 5591 9575 6452 9595
rect 4295 9539 6452 9575
rect 6508 9539 7380 9595
rect 4295 9525 7380 9539
rect -289 9377 7380 9525
rect -289 9363 6452 9377
rect -289 9307 3963 9363
rect 4019 9307 4239 9363
rect 4295 9321 6452 9363
rect 6508 9321 7380 9377
rect 4295 9307 7380 9321
rect -289 9194 7380 9307
rect -289 8151 7380 9060
rect -289 5090 7380 7813
rect 414 2234 7380 2916
rect 414 1078 7380 1986
rect 414 -1 7380 907
use M1_NACTIVE4310590878124_256x8m81  M1_NACTIVE4310590878124_256x8m81_0
timestamp 1666464484
transform 1 0 3990 0 1 9680
box 0 0 1 1
use M1_NACTIVE4310590878124_256x8m81  M1_NACTIVE4310590878124_256x8m81_1
timestamp 1666464484
transform 1 0 6482 0 1 9680
box 0 0 1 1
use M1_PACTIVE$$47509548_256x8m81  M1_PACTIVE$$47509548_256x8m81_0
timestamp 1666464484
transform 1 0 5481 0 1 11376
box -1975 -80 1975 80
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_0
timestamp 1666464484
transform 1 0 3314 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_1
timestamp 1666464484
transform 1 0 1522 0 1 3759
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_2
timestamp 1666464484
transform 1 0 2062 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_3
timestamp 1666464484
transform 1 0 3090 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_4
timestamp 1666464484
transform 1 0 494 0 1 3351
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_5
timestamp 1666464484
transform 1 0 1298 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_6
timestamp 1666464484
transform 1 0 270 0 1 3759
box 0 0 1 1
use M1_POLY2$$44753964_256x8m81  M1_POLY2$$44753964_256x8m81_7
timestamp 1666464484
transform 1 0 2286 0 1 3351
box 0 0 1 1
use M1_POLY24310590878126_256x8m81  M1_POLY24310590878126_256x8m81_0
timestamp 1666464484
transform 1 0 5985 0 1 9417
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1666464484
transform 0 -1 4242 1 0 10079
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_1
timestamp 1666464484
transform 0 -1 5170 1 0 9970
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_2
timestamp 1666464484
transform 1 0 4928 0 1 10375
box 0 0 1 1
use M2_M1$$34864172_256x8m81  M2_M1$$34864172_256x8m81_0
timestamp 1666464484
transform 1 0 5455 0 1 9367
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1666464484
transform 1 0 7122 0 1 9979
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1666464484
transform 1 0 4267 0 1 9662
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1666464484
transform 1 0 6480 0 1 9676
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1666464484
transform 1 0 3991 0 1 9662
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1666464484
transform 1 0 4926 0 1 10469
box 0 0 1 1
use M2_M1$$43375660_R90_256x8m81  M2_M1$$43375660_R90_256x8m81_0
timestamp 1666464484
transform 0 -1 5457 1 0 9603
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_0
timestamp 1666464484
transform 1 0 4267 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_1
timestamp 1666464484
transform 1 0 4706 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_256x8m81  M2_M1$$43380780_256x8m81_2
timestamp 1666464484
transform 1 0 6090 0 1 10519
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_0
timestamp 1666464484
transform 1 0 5169 0 1 3555
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_1
timestamp 1666464484
transform 1 0 6346 0 1 3353
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_2
timestamp 1666464484
transform 1 0 6860 0 1 3151
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_0
timestamp 1666464484
transform 1 0 4233 0 1 10076
box 0 0 1 1
use M2_M1431059087810_256x8m81  M2_M1431059087810_256x8m81_1
timestamp 1666464484
transform 1 0 5161 0 1 10076
box 0 0 1 1
use M3_M2$$43368492_R90_256x8m81  M3_M2$$43368492_R90_256x8m81_0
timestamp 1666464484
transform 0 -1 5457 1 0 9603
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_0
timestamp 1666464484
transform 1 0 4267 0 1 9553
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_1
timestamp 1666464484
transform 1 0 6480 0 1 9567
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_2
timestamp 1666464484
transform 1 0 4267 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_3
timestamp 1666464484
transform 1 0 4706 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_4
timestamp 1666464484
transform 1 0 3991 0 1 9553
box 0 0 1 1
use M3_M2$$47108140_256x8m81  M3_M2$$47108140_256x8m81_5
timestamp 1666464484
transform 1 0 6090 0 1 10519
box 0 0 1 1
use nmos_1p2$$46563372_256x8m81  nmos_1p2$$46563372_256x8m81_0
timestamp 1666464484
transform 1 0 5951 0 1 10236
box -119 -74 177 264
use nmos_5p04310590878140_256x8m81  nmos_5p04310590878140_256x8m81_0
timestamp 1666464484
transform 1 0 4326 0 1 10240
box -88 -44 208 318
use nmos_5p04310590878140_256x8m81  nmos_5p04310590878140_256x8m81_1
timestamp 1666464484
transform 1 0 4550 0 1 10240
box -88 -44 208 318
use pmos_5p04310590878173_256x8m81  pmos_5p04310590878173_256x8m81_0
timestamp 1666464484
transform 1 0 5802 0 1 9519
box -208 -120 552 348
use xpredec0_bot_256x8m81  xpredec0_bot_256x8m81_0
timestamp 1666464484
transform 1 0 5424 0 1 632
box -106 -633 1824 8575
use xpredec0_bot_256x8m81  xpredec0_bot_256x8m81_1
timestamp 1666464484
transform 1 0 3733 0 1 632
box -106 -633 1824 8575
use xpredec0_xa_256x8m81  xpredec0_xa_256x8m81_0
timestamp 1666464484
transform -1 0 4025 0 1 34
box 153 -35 1633 11401
use xpredec0_xa_256x8m81  xpredec0_xa_256x8m81_1
timestamp 1666464484
transform -1 0 2233 0 1 34
box 153 -35 1633 11401
use xpredec0_xa_256x8m81  xpredec0_xa_256x8m81_2
timestamp 1666464484
transform 1 0 1351 0 1 34
box 153 -35 1633 11401
use xpredec0_xa_256x8m81  xpredec0_xa_256x8m81_3
timestamp 1666464484
transform 1 0 -441 0 1 34
box 153 -35 1633 11401
<< labels >>
rlabel metal3 s 7240 9508 7240 9508 4 vdd
port 1 nsew
rlabel metal3 s 7240 10455 7240 10455 4 vss
port 2 nsew
rlabel metal3 s 7240 6422 7240 6422 4 vdd
port 1 nsew
rlabel metal3 s 7240 413 7240 413 4 vss
port 2 nsew
rlabel metal3 s 7240 1517 7240 1517 4 vdd
port 1 nsew
rlabel metal3 s 7240 2550 7240 2550 4 vss
port 2 nsew
rlabel metal3 s 7240 8587 7240 8587 4 vss
port 2 nsew
rlabel metal2 s 6911 279 6911 279 4 A[0]
port 3 nsew
rlabel metal2 s 4078 10093 4078 10093 4 men
port 4 nsew
rlabel metal2 s 2866 11124 2866 11124 4 x[0]
port 5 nsew
rlabel metal2 s 2503 11124 2503 11124 4 x[1]
port 6 nsew
rlabel metal2 s 1074 11124 1074 11124 4 x[2]
port 7 nsew
rlabel metal2 s 718 11124 718 11124 4 x[3]
port 8 nsew
rlabel metal2 s 5220 279 5220 279 4 A[1]
port 9 nsew
rlabel metal2 s 4926 10573 4926 10573 4 clk
port 10 nsew
<< properties >>
string GDS_END 1059642
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1052150
<< end >>
