magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 488 1986 1630 2449
rect 4 797 359 1986
rect 487 797 1630 1986
<< psubdiff >>
rect 149 2775 466 2834
rect 149 2729 205 2775
rect 251 2729 363 2775
rect 409 2729 466 2775
rect 149 2669 466 2729
rect 110 508 243 567
rect 110 462 153 508
rect 199 462 243 508
rect 110 345 243 462
rect 110 299 153 345
rect 199 299 243 345
rect 110 239 243 299
<< nsubdiff >>
rect 110 1801 243 1846
rect 110 1755 153 1801
rect 199 1755 243 1801
rect 110 1608 243 1755
rect 110 1562 153 1608
rect 199 1562 243 1608
rect 110 1415 243 1562
rect 110 1369 153 1415
rect 199 1369 243 1415
rect 110 1223 243 1369
rect 110 1177 153 1223
rect 199 1177 243 1223
rect 110 1015 243 1177
<< psubdiffcont >>
rect 205 2729 251 2775
rect 363 2729 409 2775
rect 153 462 199 508
rect 153 299 199 345
<< nsubdiffcont >>
rect 153 1755 199 1801
rect 153 1562 199 1608
rect 153 1369 199 1415
rect 153 1177 199 1223
<< polysilicon >>
rect 742 2339 862 2558
rect 1256 2527 1376 2588
rect 1582 2527 1666 2528
rect 1256 2509 1666 2527
rect 1256 2461 1601 2509
rect 1582 2369 1601 2461
rect 1647 2369 1666 2509
rect 375 2091 459 2110
rect 375 2045 394 2091
rect 440 2056 459 2091
rect 742 2056 862 2127
rect 440 2045 862 2056
rect 375 1996 862 2045
rect 1256 2028 1376 2087
rect 1256 2009 1439 2028
rect 1256 1963 1374 2009
rect 1420 1963 1439 2009
rect 1256 1944 1439 1963
rect 1582 1762 1666 2369
rect 1256 1693 1666 1762
rect 1256 1663 1376 1693
rect 518 864 638 908
rect 742 864 862 908
rect 518 819 1024 864
rect 518 773 904 819
rect 950 773 1024 819
rect 1490 835 1683 880
rect 1490 804 1563 835
rect 1489 803 1563 804
rect 518 727 1024 773
rect 1256 789 1563 803
rect 1609 789 1683 835
rect 1256 743 1683 789
rect 518 688 638 727
rect 742 688 862 727
rect 1256 656 1376 743
<< polycontact >>
rect 1601 2369 1647 2509
rect 394 2045 440 2091
rect 1374 1963 1420 2009
rect 904 773 950 819
rect 1563 789 1609 835
<< metal1 >>
rect 632 2864 1472 2968
rect 158 2775 457 2825
rect 158 2771 205 2775
rect 113 2731 205 2771
rect 113 2679 150 2731
rect 202 2729 205 2731
rect 251 2729 363 2775
rect 409 2729 457 2775
rect 202 2679 457 2729
rect 113 2678 457 2679
rect 113 2513 240 2678
rect 113 2461 150 2513
rect 202 2461 240 2513
rect 113 2420 240 2461
rect 632 2116 748 2864
rect 851 2731 978 2771
rect 851 2679 888 2731
rect 940 2679 978 2731
rect 851 2513 978 2679
rect 851 2461 888 2513
rect 940 2461 978 2513
rect 851 2420 978 2461
rect 383 2091 451 2102
rect 383 2045 394 2091
rect 440 2045 451 2091
rect 383 2039 451 2045
rect 359 2038 480 2039
rect 359 1946 748 2038
rect 119 1801 524 1837
rect 119 1755 153 1801
rect 199 1772 524 1801
rect 119 1720 156 1755
rect 208 1720 524 1772
rect 119 1608 524 1720
rect 119 1562 153 1608
rect 199 1562 524 1608
rect 119 1554 524 1562
rect 119 1502 156 1554
rect 208 1502 524 1554
rect 119 1415 524 1502
rect 119 1369 153 1415
rect 199 1369 524 1415
rect 119 1336 524 1369
rect 119 1284 156 1336
rect 208 1284 524 1336
rect 119 1223 524 1284
rect 119 1177 153 1223
rect 199 1177 524 1223
rect 119 947 524 1177
rect 115 609 524 649
rect 115 557 152 609
rect 204 557 524 609
rect 115 508 524 557
rect 632 539 748 1946
rect 856 1916 972 2308
rect 850 1876 978 1916
rect 850 1824 888 1876
rect 940 1824 978 1876
rect 850 1658 978 1824
rect 850 1606 888 1658
rect 940 1606 978 1658
rect 850 1440 978 1606
rect 850 1388 888 1440
rect 940 1388 978 1440
rect 850 1222 978 1388
rect 850 1170 888 1222
rect 940 1170 978 1222
rect 850 1130 978 1170
rect 1146 855 1262 2628
rect 1370 2116 1472 2864
rect 1564 2558 1691 2598
rect 1564 2369 1601 2558
rect 1653 2506 1691 2558
rect 1647 2369 1691 2506
rect 1564 2340 1691 2369
rect 1564 2288 1601 2340
rect 1653 2288 1691 2340
rect 1564 2247 1691 2288
rect 1340 2009 1691 2045
rect 1340 1963 1374 2009
rect 1420 2005 1691 2009
rect 1420 1963 1601 2005
rect 1340 1953 1601 1963
rect 1653 1953 1691 2005
rect 1340 1926 1691 1953
rect 1564 1787 1691 1926
rect 1564 1735 1601 1787
rect 1653 1735 1691 1787
rect 1564 1694 1691 1735
rect 870 819 1262 855
rect 870 773 904 819
rect 950 773 1262 819
rect 870 736 1262 773
rect 1145 735 1262 736
rect 851 609 978 649
rect 851 557 888 609
rect 940 557 978 609
rect 1146 561 1262 735
rect 1340 563 1450 1633
rect 1564 871 1644 1694
rect 1529 835 1644 871
rect 1529 789 1563 835
rect 1609 789 1644 835
rect 1529 752 1644 789
rect 115 462 153 508
rect 199 462 524 508
rect 115 391 524 462
rect 115 339 152 391
rect 204 339 524 391
rect 632 353 748 473
rect 851 391 978 557
rect 115 299 153 339
rect 199 303 524 339
rect 851 339 888 391
rect 940 339 978 391
rect 199 299 242 303
rect 115 298 242 299
rect 851 298 978 339
rect 1340 523 1485 563
rect 1340 471 1395 523
rect 1447 471 1485 523
rect 1340 305 1485 471
rect 119 248 234 298
rect 1340 253 1395 305
rect 1447 253 1485 305
rect 1340 212 1485 253
<< via1 >>
rect 150 2679 202 2731
rect 150 2461 202 2513
rect 888 2679 940 2731
rect 888 2461 940 2513
rect 156 1755 199 1772
rect 199 1755 208 1772
rect 156 1720 208 1755
rect 156 1502 208 1554
rect 156 1284 208 1336
rect 152 557 204 609
rect 888 1824 940 1876
rect 888 1606 940 1658
rect 888 1388 940 1440
rect 888 1170 940 1222
rect 1601 2509 1653 2558
rect 1601 2506 1647 2509
rect 1647 2506 1653 2509
rect 1601 2288 1653 2340
rect 1601 1953 1653 2005
rect 1601 1735 1653 1787
rect 888 557 940 609
rect 152 345 204 391
rect 152 339 153 345
rect 153 339 199 345
rect 199 339 204 345
rect 888 339 940 391
rect 1395 471 1447 523
rect 1395 253 1447 305
<< metal2 >>
rect 113 2842 240 2880
rect 113 2786 148 2842
rect 204 2786 240 2842
rect 113 2731 240 2786
rect 113 2679 150 2731
rect 202 2679 240 2731
rect 113 2624 240 2679
rect 113 2568 148 2624
rect 204 2568 240 2624
rect 113 2513 240 2568
rect 113 2461 150 2513
rect 202 2461 240 2513
rect 113 2406 240 2461
rect 113 2350 148 2406
rect 204 2350 240 2406
rect 113 2312 240 2350
rect 851 2842 978 2880
rect 851 2786 886 2842
rect 942 2786 978 2842
rect 851 2731 978 2786
rect 851 2679 888 2731
rect 940 2679 978 2731
rect 851 2624 978 2679
rect 851 2568 886 2624
rect 942 2568 978 2624
rect 851 2513 978 2568
rect 851 2461 888 2513
rect 940 2461 978 2513
rect 851 2406 978 2461
rect 851 2350 886 2406
rect 942 2350 978 2406
rect 851 2312 978 2350
rect 1564 2558 1691 2598
rect 1564 2506 1601 2558
rect 1653 2506 1691 2558
rect 1564 2340 1691 2506
rect 1564 2288 1601 2340
rect 1653 2288 1691 2340
rect 1564 2247 1691 2288
rect 1564 2005 1691 2045
rect 1564 1953 1601 2005
rect 1653 1953 1691 2005
rect 850 1878 978 1916
rect 850 1822 886 1878
rect 942 1822 978 1878
rect 119 1774 247 1812
rect 119 1718 154 1774
rect 210 1718 247 1774
rect 119 1556 247 1718
rect 119 1500 154 1556
rect 210 1500 247 1556
rect 119 1338 247 1500
rect 119 1282 154 1338
rect 210 1282 247 1338
rect 119 1244 247 1282
rect 850 1660 978 1822
rect 1564 1787 1691 1953
rect 1564 1735 1601 1787
rect 1653 1735 1691 1787
rect 1564 1694 1691 1735
rect 850 1604 886 1660
rect 942 1604 978 1660
rect 850 1442 978 1604
rect 850 1386 886 1442
rect 942 1386 978 1442
rect 850 1224 978 1386
rect 850 1168 886 1224
rect 942 1168 978 1224
rect 850 1130 978 1168
rect 114 611 242 649
rect 114 555 150 611
rect 206 555 242 611
rect 114 393 242 555
rect 114 337 150 393
rect 206 337 242 393
rect 114 298 242 337
rect 850 611 978 649
rect 850 555 886 611
rect 942 555 978 611
rect 850 393 978 555
rect 850 337 886 393
rect 942 337 978 393
rect 850 298 978 337
rect 1358 523 1485 563
rect 1358 471 1395 523
rect 1447 471 1485 523
rect 1358 305 1485 471
rect 1358 253 1395 305
rect 1447 253 1485 305
rect 1358 212 1485 253
<< via2 >>
rect 148 2786 204 2842
rect 148 2568 204 2624
rect 148 2350 204 2406
rect 886 2786 942 2842
rect 886 2568 942 2624
rect 886 2350 942 2406
rect 886 1876 942 1878
rect 886 1824 888 1876
rect 888 1824 940 1876
rect 940 1824 942 1876
rect 886 1822 942 1824
rect 154 1772 210 1774
rect 154 1720 156 1772
rect 156 1720 208 1772
rect 208 1720 210 1772
rect 154 1718 210 1720
rect 154 1554 210 1556
rect 154 1502 156 1554
rect 156 1502 208 1554
rect 208 1502 210 1554
rect 154 1500 210 1502
rect 154 1336 210 1338
rect 154 1284 156 1336
rect 156 1284 208 1336
rect 208 1284 210 1336
rect 154 1282 210 1284
rect 886 1658 942 1660
rect 886 1606 888 1658
rect 888 1606 940 1658
rect 940 1606 942 1658
rect 886 1604 942 1606
rect 886 1440 942 1442
rect 886 1388 888 1440
rect 888 1388 940 1440
rect 940 1388 942 1440
rect 886 1386 942 1388
rect 886 1222 942 1224
rect 886 1170 888 1222
rect 888 1170 940 1222
rect 940 1170 942 1222
rect 886 1168 942 1170
rect 150 609 206 611
rect 150 557 152 609
rect 152 557 204 609
rect 204 557 206 609
rect 150 555 206 557
rect 150 391 206 393
rect 150 339 152 391
rect 152 339 204 391
rect 204 339 206 391
rect 150 337 206 339
rect 886 609 942 611
rect 886 557 888 609
rect 888 557 940 609
rect 940 557 942 609
rect 886 555 942 557
rect 886 391 942 393
rect 886 339 888 391
rect 888 339 940 391
rect 940 339 942 391
rect 886 337 942 339
<< metal3 >>
rect -1 2842 1692 2916
rect -1 2786 148 2842
rect 204 2786 886 2842
rect 942 2786 1692 2842
rect -1 2624 1692 2786
rect -1 2568 148 2624
rect 204 2568 886 2624
rect 942 2568 1692 2624
rect -1 2406 1692 2568
rect -1 2350 148 2406
rect 204 2350 886 2406
rect 942 2350 1692 2406
rect -1 2234 1692 2350
rect -1 1878 1692 1986
rect -1 1822 886 1878
rect 942 1822 1692 1878
rect -1 1774 1692 1822
rect -1 1718 154 1774
rect 210 1718 1692 1774
rect -1 1660 1692 1718
rect -1 1604 886 1660
rect 942 1604 1692 1660
rect -1 1556 1692 1604
rect -1 1500 154 1556
rect 210 1500 1692 1556
rect -1 1442 1692 1500
rect -1 1386 886 1442
rect 942 1386 1692 1442
rect -1 1338 1692 1386
rect -1 1282 154 1338
rect 210 1282 1692 1338
rect -1 1224 1692 1282
rect -1 1168 886 1224
rect 942 1168 1692 1224
rect -1 1078 1692 1168
rect -90 611 1692 907
rect -90 555 150 611
rect 206 555 886 611
rect 942 555 1692 611
rect -90 393 1692 555
rect -90 337 150 393
rect 206 337 886 393
rect 942 337 1692 393
rect -90 -1 1692 337
use M1_POLY2$$44753964_155_128x8m81  M1_POLY2$$44753964_155_128x8m81_0
timestamp 1666464484
transform 1 0 927 0 1 796
box 0 0 1 1
use M1_POLY2$$44753964_155_128x8m81  M1_POLY2$$44753964_155_128x8m81_1
timestamp 1666464484
transform 1 0 1586 0 1 812
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1666464484
transform 1 0 1397 0 1 1986
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1666464484
transform 1 0 417 0 1 2068
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1666464484
transform 1 0 1624 0 1 2439
box 0 0 1 1
use M1_PSUB$$45110316_128x8m81  M1_PSUB$$45110316_128x8m81_0
timestamp 1666464484
transform 1 0 307 0 1 2752
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_0
timestamp 1666464484
transform 1 0 1627 0 1 2423
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_1
timestamp 1666464484
transform 1 0 1627 0 1 1870
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_2
timestamp 1666464484
transform 1 0 1421 0 1 388
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_3
timestamp 1666464484
transform 1 0 178 0 1 474
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_4
timestamp 1666464484
transform 1 0 914 0 1 2596
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_5
timestamp 1666464484
transform 1 0 176 0 1 2596
box 0 0 1 1
use M2_M1$$43375660_154_128x8m81  M2_M1$$43375660_154_128x8m81_6
timestamp 1666464484
transform 1 0 914 0 1 474
box 0 0 1 1
use M2_M1$$43379756_153_128x8m81  M2_M1$$43379756_153_128x8m81_0
timestamp 1666464484
transform 1 0 914 0 1 1523
box 0 0 1 1
use M2_M1$$43380780_152_128x8m81  M2_M1$$43380780_152_128x8m81_0
timestamp 1666464484
transform 1 0 182 0 1 1528
box 0 0 1 1
use M3_M2$$43368492_151_128x8m81  M3_M2$$43368492_151_128x8m81_0
timestamp 1666464484
transform 1 0 914 0 1 474
box 0 0 1 1
use M3_M2$$43368492_151_128x8m81  M3_M2$$43368492_151_128x8m81_1
timestamp 1666464484
transform 1 0 178 0 1 474
box 0 0 1 1
use M3_M2$$47108140_149_128x8m81  M3_M2$$47108140_149_128x8m81_0
timestamp 1666464484
transform 1 0 182 0 1 1528
box 0 0 1 1
use M3_M2$$47108140_149_128x8m81  M3_M2$$47108140_149_128x8m81_1
timestamp 1666464484
transform 1 0 176 0 1 2596
box 0 0 1 1
use M3_M2$$47108140_149_128x8m81  M3_M2$$47108140_149_128x8m81_2
timestamp 1666464484
transform 1 0 914 0 1 2596
box 0 0 1 1
use M3_M2$$47333420_150_128x8m81  M3_M2$$47333420_150_128x8m81_0
timestamp 1666464484
transform 1 0 914 0 1 1523
box 0 0 1 1
use nmos_1p2$$46551084_157_128x8m81  nmos_1p2$$46551084_157_128x8m81_0
timestamp 1666464484
transform 1 0 1287 0 1 204
box -119 -74 177 527
use nmos_1p2$$47329324_128x8m81  nmos_1p2$$47329324_128x8m81_0
timestamp 1666464484
transform 1 0 549 0 1 295
box -119 -74 401 436
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_0
timestamp 1666464484
transform 1 0 742 0 -1 2779
box -88 -44 208 236
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_1
timestamp 1666464484
transform 1 0 1256 0 -1 2779
box -88 -44 208 236
use pmos_1p2$$46285868_160_128x8m81  pmos_1p2$$46285868_160_128x8m81_0
timestamp 1666464484
transform 1 0 1287 0 1 1179
box -286 -142 344 595
use pmos_1p2$$47330348_161_128x8m81  pmos_1p2$$47330348_161_128x8m81_0
timestamp 1666464484
transform 1 0 1287 0 -1 2308
box -286 -141 344 322
use pmos_1p2$$47330348_161_128x8m81  pmos_1p2$$47330348_161_128x8m81_1
timestamp 1666464484
transform 1 0 773 0 -1 2308
box -286 -141 344 322
use pmos_1p2$$47331372_128x8m81  pmos_1p2$$47331372_128x8m81_0
timestamp 1666464484
transform 1 0 549 0 1 939
box -286 -142 568 1048
<< labels >>
rlabel metal3 s 202 2584 202 2584 4 vss
port 1 nsew
rlabel metal3 s 132 367 132 367 4 vss
port 1 nsew
rlabel metal3 s 156 1498 156 1498 4 vdd
port 2 nsew
rlabel metal1 s 1627 2462 1627 2462 4 enb
port 3 nsew
rlabel metal1 s 1632 1789 1632 1789 4 en
port 4 nsew
rlabel metal1 s 690 413 690 413 4 ab
port 5 nsew
rlabel metal1 s 1416 413 1416 413 4 a
port 6 nsew
<< properties >>
string GDS_END 207510
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 203076
<< end >>
