magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 6583 7408 9560 8332
rect 13849 8058 15116 8348
rect 13849 7981 15441 8058
rect 10186 7417 10786 7489
rect 13850 7408 15441 7981
rect 6583 7358 8962 7408
rect 16520 7376 21087 8303
<< mvndiff >>
rect 2123 7260 2278 7648
rect 25490 7260 25646 7648
<< mvpsubdiff >>
rect 15782 8182 16254 8239
rect 15782 8136 15837 8182
rect 15883 8136 15995 8182
rect 16041 8136 16153 8182
rect 16199 8136 16254 8182
rect 15782 8079 16254 8136
<< mvnsubdiff >>
rect 13985 8182 14931 8239
rect 13985 8136 14040 8182
rect 14086 8136 14198 8182
rect 14244 8136 14356 8182
rect 14402 8136 14514 8182
rect 14560 8136 14673 8182
rect 14719 8136 14831 8182
rect 14877 8136 14931 8182
rect 13985 8079 14931 8136
<< mvpsubdiffcont >>
rect 15837 8136 15883 8182
rect 15995 8136 16041 8182
rect 16153 8136 16199 8182
<< mvnsubdiffcont >>
rect 14040 8136 14086 8182
rect 14198 8136 14244 8182
rect 14356 8136 14402 8182
rect 14514 8136 14560 8182
rect 14673 8136 14719 8182
rect 14831 8136 14877 8182
<< polysilicon >>
rect 13623 8116 13801 8135
rect 13623 8070 13642 8116
rect 13782 8070 13801 8116
rect 15364 8164 15467 8183
rect 15364 8118 15390 8164
rect 15436 8118 15467 8164
rect 13623 8051 13801 8070
rect 6556 7896 6690 8016
rect 9314 7918 9448 8023
rect 6556 7792 6659 7896
rect 6374 7672 6690 7792
rect 9314 7778 9358 7918
rect 9404 7778 9448 7918
rect 11998 7831 12082 7850
rect 11998 7792 12017 7831
rect 9314 7673 9448 7778
rect 11043 7672 11385 7792
rect 11914 7691 12017 7792
rect 12063 7691 12082 7831
rect 11914 7672 12082 7691
rect 13664 7673 13768 8051
rect 15364 7792 15467 8118
rect 18271 7906 18355 8016
rect 13915 7672 13986 7792
rect 15305 7672 15467 7792
rect 15583 7871 15667 7890
rect 15583 7731 15602 7871
rect 15648 7792 15667 7871
rect 15648 7731 15755 7792
rect 15583 7672 15755 7731
rect 16255 7672 16656 7792
rect 17975 7672 18045 7792
rect 18271 7766 18290 7906
rect 18336 7766 18355 7906
rect 18271 7672 18355 7766
rect 21010 7792 21113 8016
rect 21010 7672 21325 7792
rect 23347 7672 23417 7792
<< polycontact >>
rect 13642 8070 13782 8116
rect 15390 8118 15436 8164
rect 9358 7778 9404 7918
rect 12017 7691 12063 7831
rect 15602 7731 15648 7871
rect 18290 7766 18336 7906
<< metal1 >>
rect 2123 7516 4017 8167
rect 4324 7852 6336 8239
rect 6728 8106 7700 8146
rect 6728 8054 6766 8106
rect 6818 8054 6977 8106
rect 7029 8054 7188 8106
rect 7240 8054 7399 8106
rect 7451 8054 7610 8106
rect 7662 8054 7700 8106
rect 6728 8014 7700 8054
rect 11385 8131 11913 8219
rect 11385 8079 11575 8131
rect 11627 8079 11755 8131
rect 11807 8079 11913 8131
rect 9323 7918 9439 7985
rect 6482 7788 6767 7908
rect 4335 7645 5307 7685
rect 6482 7677 6598 7788
rect 9323 7778 9358 7918
rect 9404 7778 9439 7918
rect 10338 7908 10888 7915
rect 10337 7874 10888 7908
rect 10337 7822 10376 7874
rect 10428 7822 10587 7874
rect 10639 7822 10798 7874
rect 10850 7822 10888 7874
rect 10337 7788 10888 7822
rect 11385 7913 11913 8079
rect 13531 8182 14912 8219
rect 15755 8218 16283 8219
rect 13531 8178 14040 8182
rect 13531 8126 14033 8178
rect 14086 8136 14198 8182
rect 14244 8178 14356 8182
rect 14085 8126 14244 8136
rect 14296 8136 14356 8178
rect 14402 8178 14514 8182
rect 14402 8136 14455 8178
rect 14296 8126 14455 8136
rect 14507 8136 14514 8178
rect 14560 8136 14673 8182
rect 14719 8136 14831 8182
rect 14877 8136 14912 8182
rect 14507 8126 14912 8136
rect 13531 8117 14912 8126
rect 13531 8065 13569 8117
rect 13621 8116 13781 8117
rect 13621 8070 13642 8116
rect 13833 8099 14912 8117
rect 15061 8182 16283 8218
rect 15061 8178 15837 8182
rect 15061 8126 15100 8178
rect 15152 8126 15311 8178
rect 15363 8164 15522 8178
rect 15363 8126 15390 8164
rect 15061 8118 15390 8126
rect 15436 8126 15522 8164
rect 15574 8126 15733 8178
rect 15785 8136 15837 8178
rect 15883 8136 15995 8182
rect 16041 8136 16153 8182
rect 16199 8136 16283 8182
rect 20112 8140 20874 8146
rect 15785 8126 16283 8136
rect 15436 8118 16283 8126
rect 13833 8086 14545 8099
rect 13833 8085 14040 8086
rect 15061 8085 16283 8118
rect 13621 8065 13781 8070
rect 13833 8065 13871 8085
rect 13531 8024 13871 8065
rect 11385 7861 11575 7913
rect 11627 7861 11755 7913
rect 11807 7861 11913 7913
rect 15591 7871 15659 7882
rect 11385 7821 11913 7861
rect 12006 7831 12334 7868
rect 10338 7782 10888 7788
rect 4335 7593 4373 7645
rect 4425 7593 4584 7645
rect 4636 7593 4795 7645
rect 4847 7593 5006 7645
rect 5058 7593 5217 7645
rect 5269 7593 5307 7645
rect 4335 7553 5307 7593
rect 6240 7557 6598 7677
rect 6728 7643 7700 7683
rect 6728 7591 6766 7643
rect 6818 7591 6977 7643
rect 7029 7591 7188 7643
rect 7240 7591 7399 7643
rect 7451 7591 7610 7643
rect 7662 7591 7700 7643
rect 6728 7551 7700 7591
rect 9323 7677 9439 7778
rect 12006 7691 12017 7831
rect 12063 7822 12334 7831
rect 13509 7822 14174 7868
rect 15591 7867 15602 7871
rect 12063 7691 12074 7822
rect 15268 7821 15602 7867
rect 15591 7731 15602 7821
rect 15648 7731 15659 7871
rect 15755 7788 16283 8085
rect 16656 8106 20942 8140
rect 16656 8054 20151 8106
rect 20203 8054 20362 8106
rect 20414 8054 20573 8106
rect 20625 8054 20784 8106
rect 20836 8054 20942 8106
rect 16656 8020 20942 8054
rect 16656 7836 17974 8020
rect 20112 8013 20874 8020
rect 18279 7906 18347 7917
rect 15591 7720 15659 7731
rect 18279 7766 18290 7906
rect 18336 7766 18347 7906
rect 20898 7821 21184 7867
rect 18279 7755 18347 7766
rect 12006 7680 12074 7691
rect 9323 7557 11913 7677
rect 12294 7643 13478 7684
rect 18279 7677 18346 7755
rect 12294 7591 12333 7643
rect 12385 7591 12544 7643
rect 12596 7591 12755 7643
rect 12807 7591 12966 7643
rect 13018 7591 13177 7643
rect 13229 7591 13387 7643
rect 13439 7591 13478 7643
rect 13570 7598 14174 7644
rect 12294 7550 13478 7591
rect 15755 7557 18346 7677
rect 20112 7643 20874 7683
rect 20112 7591 20151 7643
rect 20203 7591 20362 7643
rect 20414 7591 20573 7643
rect 20625 7591 20784 7643
rect 20836 7591 20874 7643
rect 21067 7643 21184 7821
rect 21324 7802 23346 8219
rect 22366 7643 23338 7683
rect 21067 7597 21425 7643
rect 20112 7550 20874 7591
rect 22366 7591 22404 7643
rect 22456 7591 22615 7643
rect 22667 7591 22826 7643
rect 22878 7591 23037 7643
rect 23089 7591 23248 7643
rect 23300 7591 23338 7643
rect 22366 7551 23338 7591
rect 23751 7516 25646 8167
rect 2123 7265 2278 7516
rect 25490 7265 25646 7516
rect 13220 6988 13349 7028
rect 13220 6936 13258 6988
rect 13310 6936 13349 6988
rect 13220 6909 13349 6936
rect 13220 6896 13348 6909
rect 14730 6757 14859 6797
rect 14730 6705 14768 6757
rect 14820 6705 14859 6757
rect 14730 6678 14859 6705
rect 14730 6665 14858 6678
rect 16882 6648 17011 6688
rect 16882 6596 16920 6648
rect 16972 6596 17011 6648
rect 16882 6569 17011 6596
rect 16882 6556 17010 6569
rect 17260 6004 17389 6044
rect 17260 5952 17298 6004
rect 17350 5952 17389 6004
rect 14730 5895 14859 5935
rect 17260 5925 17389 5952
rect 17260 5912 17388 5925
rect 14730 5843 14768 5895
rect 14820 5843 14859 5895
rect 14730 5816 14859 5843
rect 14730 5803 14858 5816
rect 13220 5664 13349 5704
rect 13220 5612 13258 5664
rect 13310 5612 13349 5664
rect 13220 5585 13349 5612
rect 13220 5572 13348 5585
rect 13220 5188 13349 5228
rect 13220 5136 13258 5188
rect 13310 5136 13349 5188
rect 13220 5109 13349 5136
rect 13220 5096 13348 5109
rect 14730 4957 14859 4997
rect 14730 4905 14768 4957
rect 14820 4905 14859 4957
rect 14730 4878 14859 4905
rect 14730 4865 14858 4878
rect 17638 4848 17767 4888
rect 17638 4796 17676 4848
rect 17728 4796 17767 4848
rect 17638 4769 17767 4796
rect 17638 4756 17766 4769
rect 18016 4204 18145 4244
rect 18016 4152 18054 4204
rect 18106 4152 18145 4204
rect 14730 4095 14859 4135
rect 18016 4125 18145 4152
rect 18016 4112 18144 4125
rect 14730 4043 14768 4095
rect 14820 4043 14859 4095
rect 14730 4016 14859 4043
rect 14730 4003 14858 4016
rect 13220 3864 13349 3904
rect 13220 3812 13258 3864
rect 13310 3812 13349 3864
rect 13220 3785 13349 3812
rect 13220 3772 13348 3785
rect 13220 3388 13349 3428
rect 13220 3336 13258 3388
rect 13310 3336 13349 3388
rect 13220 3309 13349 3336
rect 13220 3296 13348 3309
rect 14730 3157 14859 3197
rect 14730 3105 14768 3157
rect 14820 3105 14859 3157
rect 14730 3078 14859 3105
rect 14730 3065 14858 3078
rect 18393 3048 18522 3088
rect 18393 2996 18431 3048
rect 18483 2996 18522 3048
rect 18393 2969 18522 2996
rect 18393 2956 18521 2969
rect 18771 2404 18900 2444
rect 18771 2352 18809 2404
rect 18861 2352 18900 2404
rect 14730 2295 14859 2335
rect 18771 2325 18900 2352
rect 18771 2312 18899 2325
rect 14730 2243 14768 2295
rect 14820 2243 14859 2295
rect 14730 2216 14859 2243
rect 14730 2203 14858 2216
rect 13220 2064 13349 2104
rect 13220 2012 13258 2064
rect 13310 2012 13349 2064
rect 13220 1985 13349 2012
rect 13220 1972 13348 1985
rect 13220 1588 13349 1628
rect 13220 1536 13258 1588
rect 13310 1536 13349 1588
rect 13220 1509 13349 1536
rect 13220 1496 13348 1509
rect 14730 1357 14859 1397
rect 14730 1305 14768 1357
rect 14820 1305 14859 1357
rect 14730 1278 14859 1305
rect 14730 1265 14858 1278
rect 19149 1248 19278 1288
rect 19149 1196 19187 1248
rect 19239 1196 19278 1248
rect 19149 1169 19278 1196
rect 19149 1156 19277 1169
rect 19526 604 19655 644
rect 19526 552 19564 604
rect 19616 552 19655 604
rect 14730 495 14859 535
rect 19526 525 19655 552
rect 19526 512 19654 525
rect 14730 443 14768 495
rect 14820 443 14859 495
rect 14730 416 14859 443
rect 14730 403 14858 416
rect 13220 264 13349 304
rect 13220 212 13258 264
rect 13310 212 13349 264
rect 13220 185 13349 212
rect 13220 172 13348 185
<< via1 >>
rect 6766 8054 6818 8106
rect 6977 8054 7029 8106
rect 7188 8054 7240 8106
rect 7399 8054 7451 8106
rect 7610 8054 7662 8106
rect 11575 8079 11627 8131
rect 11755 8079 11807 8131
rect 10376 7822 10428 7874
rect 10587 7822 10639 7874
rect 10798 7822 10850 7874
rect 14033 8136 14040 8178
rect 14040 8136 14085 8178
rect 14033 8126 14085 8136
rect 14244 8126 14296 8178
rect 14455 8126 14507 8178
rect 13569 8065 13621 8117
rect 13781 8116 13833 8117
rect 13781 8070 13782 8116
rect 13782 8070 13833 8116
rect 15100 8126 15152 8178
rect 15311 8126 15363 8178
rect 15522 8126 15574 8178
rect 15733 8126 15785 8178
rect 13781 8065 13833 8070
rect 11575 7861 11627 7913
rect 11755 7861 11807 7913
rect 4373 7593 4425 7645
rect 4584 7593 4636 7645
rect 4795 7593 4847 7645
rect 5006 7593 5058 7645
rect 5217 7593 5269 7645
rect 6766 7591 6818 7643
rect 6977 7591 7029 7643
rect 7188 7591 7240 7643
rect 7399 7591 7451 7643
rect 7610 7591 7662 7643
rect 20151 8054 20203 8106
rect 20362 8054 20414 8106
rect 20573 8054 20625 8106
rect 20784 8054 20836 8106
rect 12333 7591 12385 7643
rect 12544 7591 12596 7643
rect 12755 7591 12807 7643
rect 12966 7591 13018 7643
rect 13177 7591 13229 7643
rect 13387 7591 13439 7643
rect 20151 7591 20203 7643
rect 20362 7591 20414 7643
rect 20573 7591 20625 7643
rect 20784 7591 20836 7643
rect 22404 7591 22456 7643
rect 22615 7591 22667 7643
rect 22826 7591 22878 7643
rect 23037 7591 23089 7643
rect 23248 7591 23300 7643
rect 13258 6936 13310 6988
rect 14768 6705 14820 6757
rect 16920 6596 16972 6648
rect 17298 5952 17350 6004
rect 14768 5843 14820 5895
rect 13258 5612 13310 5664
rect 13258 5136 13310 5188
rect 14768 4905 14820 4957
rect 17676 4796 17728 4848
rect 18054 4152 18106 4204
rect 14768 4043 14820 4095
rect 13258 3812 13310 3864
rect 13258 3336 13310 3388
rect 14768 3105 14820 3157
rect 18431 2996 18483 3048
rect 18809 2352 18861 2404
rect 14768 2243 14820 2295
rect 13258 2012 13310 2064
rect 13258 1536 13310 1588
rect 14768 1305 14820 1357
rect 19187 1196 19239 1248
rect 19564 552 19616 604
rect 14768 443 14820 495
rect 13258 212 13310 264
<< metal2 >>
rect 2092 7213 4211 8276
rect 5550 8128 6347 8201
rect 5550 8072 5611 8128
rect 5667 8072 5822 8128
rect 5878 8072 6033 8128
rect 6089 8072 6244 8128
rect 6300 8072 6347 8128
rect 4334 7647 5307 7686
rect 4334 7591 4371 7647
rect 4427 7591 4582 7647
rect 4638 7591 4793 7647
rect 4849 7591 5004 7647
rect 5060 7591 5215 7647
rect 5271 7591 5307 7647
rect 4334 7553 5307 7591
rect 5550 7213 6347 8072
rect 6451 8106 7738 8201
rect 6451 8054 6766 8106
rect 6818 8054 6977 8106
rect 7029 8054 7188 8106
rect 7240 8054 7399 8106
rect 7451 8054 7610 8106
rect 7662 8054 7738 8106
rect 6451 7643 7738 8054
rect 6451 7591 6766 7643
rect 6818 7591 6977 7643
rect 7029 7591 7188 7643
rect 7240 7591 7399 7643
rect 7451 7591 7610 7643
rect 7662 7591 7738 7643
rect 6451 7213 7738 7591
rect 8186 7645 9066 7684
rect 8186 7589 8222 7645
rect 8278 7589 8433 7645
rect 8489 7589 8644 7645
rect 8700 7589 8855 7645
rect 8911 7589 9066 7645
rect 8186 7213 9066 7589
rect 9591 7213 10186 8201
rect 10276 7874 10941 8201
rect 10276 7822 10376 7874
rect 10428 7822 10587 7874
rect 10639 7822 10798 7874
rect 10850 7822 10941 7874
rect 10276 7213 10941 7822
rect 11537 8131 11846 8201
rect 13994 8178 14545 8219
rect 11537 8128 11575 8131
rect 11627 8128 11755 8131
rect 11807 8128 11846 8131
rect 11537 8072 11573 8128
rect 11629 8072 11753 8128
rect 11809 8072 11846 8128
rect 11537 7913 11846 8072
rect 13531 8117 13871 8158
rect 13531 8065 13569 8117
rect 13621 8065 13781 8117
rect 13833 8065 13871 8117
rect 13531 8024 13871 8065
rect 13994 8126 14033 8178
rect 14085 8126 14244 8178
rect 14296 8126 14455 8178
rect 14507 8126 14545 8178
rect 11537 7861 11575 7913
rect 11627 7861 11755 7913
rect 11807 7861 11846 7913
rect 11537 7213 11846 7861
rect 12294 7645 13478 7684
rect 12294 7589 12331 7645
rect 12387 7589 12542 7645
rect 12598 7589 12753 7645
rect 12809 7589 12964 7645
rect 13020 7589 13175 7645
rect 13231 7589 13385 7645
rect 13441 7589 13478 7645
rect 12294 7550 13478 7589
rect 13994 7638 14545 8126
rect 13994 7582 14031 7638
rect 14087 7582 14242 7638
rect 14298 7582 14453 7638
rect 14509 7582 14545 7638
rect 13994 7364 14545 7582
rect 15026 8178 15887 8219
rect 15026 8126 15100 8178
rect 15152 8126 15311 8178
rect 15363 8126 15522 8178
rect 15574 8126 15733 8178
rect 15785 8126 15887 8178
rect 12040 7228 12639 7364
rect 12040 7172 12100 7228
rect 12156 7172 12311 7228
rect 12367 7172 12522 7228
rect 12578 7172 12639 7228
rect 12040 7099 12639 7172
rect 12880 7123 14823 7364
rect 15026 7213 15887 8126
rect 20112 8106 21313 8201
rect 20112 8054 20151 8106
rect 20203 8054 20362 8106
rect 20414 8054 20573 8106
rect 20625 8054 20784 8106
rect 20836 8054 21313 8106
rect 20112 7643 21313 8054
rect 20112 7591 20151 7643
rect 20203 7591 20362 7643
rect 20414 7591 20573 7643
rect 20625 7591 20784 7643
rect 20836 7591 21313 7643
rect 20112 7213 21313 7591
rect 21421 8128 22236 8219
rect 21421 8072 21458 8128
rect 21514 8072 21669 8128
rect 21725 8072 21880 8128
rect 21936 8072 22091 8128
rect 22147 8072 22236 8128
rect 21421 7213 22236 8072
rect 22365 7645 23338 7684
rect 22365 7589 22402 7645
rect 22458 7589 22613 7645
rect 22669 7589 22824 7645
rect 22880 7589 23035 7645
rect 23091 7589 23246 7645
rect 23302 7589 23338 7645
rect 22365 7551 23338 7589
rect 23549 7213 25677 8276
rect 13220 6988 13348 7029
rect 13220 6936 13258 6988
rect 13310 6936 13348 6988
rect 13220 6895 13348 6936
rect 14730 6757 14858 6798
rect 14730 6705 14768 6757
rect 14820 6705 14858 6757
rect 14730 6664 14858 6705
rect 16882 6648 17010 6689
rect 16882 6596 16920 6648
rect 16972 6596 17010 6648
rect 16882 6555 17010 6596
rect 17260 6004 17388 6045
rect 17260 5952 17298 6004
rect 17350 5952 17388 6004
rect 14730 5895 14858 5936
rect 17260 5911 17388 5952
rect 14730 5843 14768 5895
rect 14820 5843 14858 5895
rect 14730 5802 14858 5843
rect 13220 5664 13348 5705
rect 13220 5612 13258 5664
rect 13310 5612 13348 5664
rect 13220 5571 13348 5612
rect 13220 5188 13348 5229
rect 13220 5136 13258 5188
rect 13310 5136 13348 5188
rect 13220 5095 13348 5136
rect 14730 4957 14858 4998
rect 14730 4905 14768 4957
rect 14820 4905 14858 4957
rect 14730 4864 14858 4905
rect 17638 4848 17766 4889
rect 17638 4796 17676 4848
rect 17728 4796 17766 4848
rect 17638 4755 17766 4796
rect 18016 4204 18144 4245
rect 18016 4152 18054 4204
rect 18106 4152 18144 4204
rect 14730 4095 14858 4136
rect 18016 4111 18144 4152
rect 14730 4043 14768 4095
rect 14820 4043 14858 4095
rect 14730 4002 14858 4043
rect 13220 3864 13348 3905
rect 13220 3812 13258 3864
rect 13310 3812 13348 3864
rect 13220 3771 13348 3812
rect 13220 3388 13348 3429
rect 13220 3336 13258 3388
rect 13310 3336 13348 3388
rect 13220 3295 13348 3336
rect 14730 3157 14858 3198
rect 14730 3105 14768 3157
rect 14820 3105 14858 3157
rect 14730 3064 14858 3105
rect 18393 3048 18521 3089
rect 18393 2996 18431 3048
rect 18483 2996 18521 3048
rect 18393 2955 18521 2996
rect 18771 2404 18899 2445
rect 18771 2352 18809 2404
rect 18861 2352 18899 2404
rect 14730 2295 14858 2336
rect 18771 2311 18899 2352
rect 14730 2243 14768 2295
rect 14820 2243 14858 2295
rect 14730 2202 14858 2243
rect 13220 2064 13348 2105
rect 13220 2012 13258 2064
rect 13310 2012 13348 2064
rect 13220 1971 13348 2012
rect 13220 1588 13348 1629
rect 13220 1536 13258 1588
rect 13310 1536 13348 1588
rect 13220 1495 13348 1536
rect 14730 1357 14858 1398
rect 14730 1305 14768 1357
rect 14820 1305 14858 1357
rect 14730 1264 14858 1305
rect 19149 1248 19277 1289
rect 19149 1196 19187 1248
rect 19239 1196 19277 1248
rect 19149 1155 19277 1196
rect 19526 604 19654 645
rect 19526 552 19564 604
rect 19616 552 19654 604
rect 14730 495 14858 536
rect 19526 511 19654 552
rect 14730 443 14768 495
rect 14820 443 14858 495
rect 14730 402 14858 443
rect 13219 264 13348 305
rect 13219 212 13258 264
rect 13310 212 13348 264
rect 13219 171 13348 212
rect 13597 171 13726 305
rect 13974 171 14104 305
rect 14352 171 14481 305
rect 14730 171 14859 305
rect 16882 171 17011 305
rect 17260 171 17389 305
rect 17637 171 17767 305
rect 18015 171 18144 305
rect 18393 171 18522 305
rect 18770 171 18900 305
rect 19148 171 19277 305
rect 19526 171 19655 305
rect 8561 -21 8691 112
rect 12841 -164 12971 -31
rect 13219 -164 13348 -31
rect 13597 -164 13726 -31
rect 13974 -164 14104 -31
rect 14352 -164 14481 -31
rect 14730 -164 14859 -31
rect 16882 -164 17011 -31
rect 17260 -164 17389 -31
rect 17637 -164 17767 -31
rect 18015 -164 18144 -31
rect 18393 -164 18522 -31
rect 18770 -164 18900 -31
rect 19148 -164 19277 -31
rect 19526 -164 19655 -31
<< via2 >>
rect 5611 8072 5667 8128
rect 5822 8072 5878 8128
rect 6033 8072 6089 8128
rect 6244 8072 6300 8128
rect 4371 7645 4427 7647
rect 4371 7593 4373 7645
rect 4373 7593 4425 7645
rect 4425 7593 4427 7645
rect 4371 7591 4427 7593
rect 4582 7645 4638 7647
rect 4582 7593 4584 7645
rect 4584 7593 4636 7645
rect 4636 7593 4638 7645
rect 4582 7591 4638 7593
rect 4793 7645 4849 7647
rect 4793 7593 4795 7645
rect 4795 7593 4847 7645
rect 4847 7593 4849 7645
rect 4793 7591 4849 7593
rect 5004 7645 5060 7647
rect 5004 7593 5006 7645
rect 5006 7593 5058 7645
rect 5058 7593 5060 7645
rect 5004 7591 5060 7593
rect 5215 7645 5271 7647
rect 5215 7593 5217 7645
rect 5217 7593 5269 7645
rect 5269 7593 5271 7645
rect 5215 7591 5271 7593
rect 8222 7589 8278 7645
rect 8433 7589 8489 7645
rect 8644 7589 8700 7645
rect 8855 7589 8911 7645
rect 11573 8079 11575 8128
rect 11575 8079 11627 8128
rect 11627 8079 11629 8128
rect 11573 8072 11629 8079
rect 11753 8079 11755 8128
rect 11755 8079 11807 8128
rect 11807 8079 11809 8128
rect 11753 8072 11809 8079
rect 12331 7643 12387 7645
rect 12331 7591 12333 7643
rect 12333 7591 12385 7643
rect 12385 7591 12387 7643
rect 12331 7589 12387 7591
rect 12542 7643 12598 7645
rect 12542 7591 12544 7643
rect 12544 7591 12596 7643
rect 12596 7591 12598 7643
rect 12542 7589 12598 7591
rect 12753 7643 12809 7645
rect 12753 7591 12755 7643
rect 12755 7591 12807 7643
rect 12807 7591 12809 7643
rect 12753 7589 12809 7591
rect 12964 7643 13020 7645
rect 12964 7591 12966 7643
rect 12966 7591 13018 7643
rect 13018 7591 13020 7643
rect 12964 7589 13020 7591
rect 13175 7643 13231 7645
rect 13175 7591 13177 7643
rect 13177 7591 13229 7643
rect 13229 7591 13231 7643
rect 13175 7589 13231 7591
rect 13385 7643 13441 7645
rect 13385 7591 13387 7643
rect 13387 7591 13439 7643
rect 13439 7591 13441 7643
rect 13385 7589 13441 7591
rect 14031 7582 14087 7638
rect 14242 7582 14298 7638
rect 14453 7582 14509 7638
rect 12100 7172 12156 7228
rect 12311 7172 12367 7228
rect 12522 7172 12578 7228
rect 21458 8072 21514 8128
rect 21669 8072 21725 8128
rect 21880 8072 21936 8128
rect 22091 8072 22147 8128
rect 22402 7643 22458 7645
rect 22402 7591 22404 7643
rect 22404 7591 22456 7643
rect 22456 7591 22458 7643
rect 22402 7589 22458 7591
rect 22613 7643 22669 7645
rect 22613 7591 22615 7643
rect 22615 7591 22667 7643
rect 22667 7591 22669 7643
rect 22613 7589 22669 7591
rect 22824 7643 22880 7645
rect 22824 7591 22826 7643
rect 22826 7591 22878 7643
rect 22878 7591 22880 7643
rect 22824 7589 22880 7591
rect 23035 7643 23091 7645
rect 23035 7591 23037 7643
rect 23037 7591 23089 7643
rect 23089 7591 23091 7643
rect 23035 7589 23091 7591
rect 23246 7643 23302 7645
rect 23246 7591 23248 7643
rect 23248 7591 23300 7643
rect 23300 7591 23302 7643
rect 23246 7589 23302 7591
<< metal3 >>
rect 69 8033 199 8167
rect 1725 8128 25945 8201
rect 1725 8072 5611 8128
rect 5667 8072 5822 8128
rect 5878 8072 6033 8128
rect 6089 8072 6244 8128
rect 6300 8072 11573 8128
rect 11629 8072 11753 8128
rect 11809 8072 21458 8128
rect 21514 8072 21669 8128
rect 21725 8072 21880 8128
rect 21936 8072 22091 8128
rect 22147 8072 25945 8128
rect 1725 7999 25945 8072
rect -1 7573 128 7707
rect 1725 7647 5307 7741
rect 1725 7591 4371 7647
rect 4427 7591 4582 7647
rect 4638 7591 4793 7647
rect 4849 7591 5004 7647
rect 5060 7591 5215 7647
rect 5271 7591 5307 7647
rect 1725 7539 5307 7591
rect 8186 7645 13478 7684
rect 8186 7589 8222 7645
rect 8278 7589 8433 7645
rect 8489 7589 8644 7645
rect 8700 7589 8855 7645
rect 8911 7589 12331 7645
rect 12387 7589 12542 7645
rect 12598 7589 12753 7645
rect 12809 7589 12964 7645
rect 13020 7589 13175 7645
rect 13231 7589 13385 7645
rect 13441 7589 13478 7645
rect 8186 7550 13478 7589
rect 13994 7638 14545 7677
rect 13994 7582 14031 7638
rect 14087 7582 14242 7638
rect 14298 7582 14453 7638
rect 14509 7582 14545 7638
rect 69 7133 199 7267
rect 12063 7228 12615 7267
rect 13994 7232 14545 7582
rect 22365 7645 25945 7741
rect 22365 7589 22402 7645
rect 22458 7589 22613 7645
rect 22669 7589 22824 7645
rect 22880 7589 23035 7645
rect 23091 7589 23246 7645
rect 23302 7589 25945 7645
rect 22365 7539 25945 7589
rect 27640 7573 27769 7707
rect 12063 7172 12100 7228
rect 12156 7172 12311 7228
rect 12367 7172 12522 7228
rect 12578 7172 12615 7228
rect 12063 7133 12615 7172
rect -1 6673 128 6807
rect 2491 6693 2621 6827
rect 25084 6693 25213 6827
rect 27640 6673 27769 6807
rect -1 5793 128 5927
rect 2491 5773 2621 5907
rect 25084 5773 25213 5907
rect 27640 5793 27769 5927
rect -1 4873 128 5007
rect 2491 4893 2621 5027
rect 25084 4893 25213 5027
rect 27640 4873 27769 5007
rect -1 3993 128 4127
rect 2491 3973 2621 4107
rect 25084 3973 25213 4107
rect 27640 3993 27769 4127
rect -1 3073 128 3207
rect 2491 3093 2621 3227
rect 25084 3093 25213 3227
rect 27640 3073 27769 3207
rect -1 2193 128 2327
rect 2491 2173 2621 2307
rect 25084 2173 25213 2307
rect 27640 2193 27769 2327
rect -1 1273 128 1407
rect 2491 1293 2621 1427
rect 25084 1293 25213 1427
rect 27640 1273 27769 1407
rect -1 393 128 527
rect 2491 373 2621 507
rect 27640 393 27769 527
use M1_NACTIVE$$203393068_64x8m81  M1_NACTIVE$$203393068_64x8m81_0
timestamp 1666464484
transform 1 0 14063 0 1 8159
box 0 0 1 1
use M1_NWELL$$204218412_64x8m81  M1_NWELL$$204218412_64x8m81_0
timestamp 1666464484
transform -1 0 25568 0 1 8086
box -221 -717 1960 228
use M1_NWELL$$204218412_64x8m81  M1_NWELL$$204218412_64x8m81_1
timestamp 1666464484
transform 1 0 2200 0 1 8086
box -221 -717 1960 228
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_0
timestamp 1666464484
transform 1 0 11463 0 1 8159
box -78 -80 1817 80
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_1
timestamp 1666464484
transform 1 0 21475 0 1 8159
box -78 -80 1817 80
use M1_PACTIVE$$204148780_64x8m81  M1_PACTIVE$$204148780_64x8m81_2
timestamp 1666464484
transform 1 0 4390 0 1 8159
box -78 -80 1817 80
use M1_PACTIVE$$204149804_64x8m81  M1_PACTIVE$$204149804_64x8m81_0
timestamp 1666464484
transform 1 0 15860 0 1 8159
box 0 0 1 1
use M1_POLY2$$204150828_64x8m81  M1_POLY2$$204150828_64x8m81_0
timestamp 1666464484
transform 1 0 9381 0 1 7848
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1666464484
transform 1 0 15413 0 1 8141
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1666464484
transform 0 -1 13712 1 0 8093
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_1
timestamp 1666464484
transform 1 0 15625 0 1 7801
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_2
timestamp 1666464484
transform 1 0 18313 0 1 7836
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_3
timestamp 1666464484
transform 1 0 12040 0 1 7761
box 0 0 1 1
use M2_M1$$201262124_64x8m81  M2_M1$$201262124_64x8m81_0
timestamp 1666464484
transform 1 0 13701 0 1 8091
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_0
timestamp 1666464484
transform 1 0 13284 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_1
timestamp 1666464484
transform 1 0 13284 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_2
timestamp 1666464484
transform 1 0 13284 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_3
timestamp 1666464484
transform 1 0 14794 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_4
timestamp 1666464484
transform 1 0 14794 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_5
timestamp 1666464484
transform 1 0 14794 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_6
timestamp 1666464484
transform 1 0 14794 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_7
timestamp 1666464484
transform 1 0 14794 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_8
timestamp 1666464484
transform 1 0 14794 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_9
timestamp 1666464484
transform 1 0 14794 0 1 469
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_10
timestamp 1666464484
transform 1 0 13284 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_11
timestamp 1666464484
transform 1 0 13284 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_12
timestamp 1666464484
transform 1 0 13284 0 1 238
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_13
timestamp 1666464484
transform 1 0 13284 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_14
timestamp 1666464484
transform 1 0 13284 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_15
timestamp 1666464484
transform 1 0 19590 0 1 578
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_16
timestamp 1666464484
transform 1 0 19213 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_17
timestamp 1666464484
transform 1 0 18835 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_18
timestamp 1666464484
transform 1 0 18457 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_19
timestamp 1666464484
transform 1 0 18080 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_20
timestamp 1666464484
transform 1 0 17702 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_21
timestamp 1666464484
transform 1 0 17324 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_22
timestamp 1666464484
transform 1 0 16946 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_23
timestamp 1666464484
transform 1 0 14794 0 1 6731
box 0 0 1 1
use M2_M1$$204138540_64x8m81  M2_M1$$204138540_64x8m81_0
timestamp 1666464484
transform 1 0 10402 0 1 7848
box 0 0 1 1
use M2_M1$$204138540_64x8m81  M2_M1$$204138540_64x8m81_1
timestamp 1666464484
transform 1 0 14059 0 1 8152
box 0 0 1 1
use M2_M1$$204139564_64x8m81  M2_M1$$204139564_64x8m81_0
timestamp 1666464484
transform 1 0 11601 0 1 8105
box 0 0 1 1
use M2_M1$$204140588_64x8m81  M2_M1$$204140588_64x8m81_0
timestamp 1666464484
transform 1 0 12359 0 1 7617
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_0
timestamp 1666464484
transform 1 0 15126 0 1 8152
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_1
timestamp 1666464484
transform 1 0 20177 0 1 8080
box 0 0 1 1
use M2_M1$$204141612_64x8m81  M2_M1$$204141612_64x8m81_2
timestamp 1666464484
transform 1 0 20177 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_0
timestamp 1666464484
transform 1 0 6792 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_1
timestamp 1666464484
transform 1 0 22430 0 1 7617
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_2
timestamp 1666464484
transform 1 0 4399 0 1 7619
box 0 0 1 1
use M2_M1$$204220460_64x8m81  M2_M1$$204220460_64x8m81_3
timestamp 1666464484
transform 1 0 6792 0 1 8080
box 0 0 1 1
use M2_M1$$204221484_64x8m81  M2_M1$$204221484_64x8m81_0
timestamp 1666464484
transform -1 0 25612 0 1 8100
box -65 -502 1751 67
use M2_M1$$204221484_64x8m81  M2_M1$$204221484_64x8m81_1
timestamp 1666464484
transform 1 0 2156 0 1 8100
box -65 -502 1751 67
use M2_M1$$204222508_64x8m81  M2_M1$$204222508_64x8m81_0
timestamp 1666464484
transform 1 0 21486 0 1 8100
box -65 -284 697 67
use M2_M1$$204222508_64x8m81  M2_M1$$204222508_64x8m81_1
timestamp 1666464484
transform 1 0 5639 0 1 8100
box -65 -284 697 67
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_0
timestamp 1666464484
transform 1 0 5639 0 1 8100
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_1
timestamp 1666464484
transform 1 0 8250 0 1 7617
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_2
timestamp 1666464484
transform 1 0 21486 0 1 8100
box 0 0 1 1
use M3_M2$$204142636_64x8m81  M3_M2$$204142636_64x8m81_3
timestamp 1666464484
transform 1 0 21486 0 1 8100
box 0 0 1 1
use M3_M2$$204143660_64x8m81  M3_M2$$204143660_64x8m81_0
timestamp 1666464484
transform 1 0 11601 0 1 8100
box 0 0 1 1
use M3_M2$$204144684_64x8m81  M3_M2$$204144684_64x8m81_0
timestamp 1666464484
transform 1 0 22430 0 1 7617
box 0 0 1 1
use M3_M2$$204144684_64x8m81  M3_M2$$204144684_64x8m81_1
timestamp 1666464484
transform 1 0 4399 0 1 7619
box 0 0 1 1
use M3_M2$$204145708_64x8m81  M3_M2$$204145708_64x8m81_0
timestamp 1666464484
transform 1 0 12359 0 1 7617
box 0 0 1 1
use M3_M2$$204146732_64x8m81  M3_M2$$204146732_64x8m81_0
timestamp 1666464484
transform 1 0 14059 0 1 7610
box 0 0 1 1
use M3_M2$$204147756_64x8m81  M3_M2$$204147756_64x8m81_0
timestamp 1666464484
transform 1 0 12339 0 1 7200
box 0 0 1 1
use nmos_1p2$$204215_R270_64x8m81  nmos_1p2$$204215_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 13604 -1 0 7762
box -119 -71 177 1389
use nmos_1p2$$204213292_R90_64x8m81  nmos_1p2$$204213292_R90_64x8m81_0
timestamp 1666464484
transform 0 -1 6346 1 0 7703
box -119 -71 177 2091
use nmos_5p04310589983299_64x8m81  nmos_5p04310589983299_64x8m81_0
timestamp 1666464484
transform 0 -1 23346 1 0 7672
box -88 -44 208 2066
use nmos_5p043105899832103_64x8m81  nmos_5p043105899832103_64x8m81_0
timestamp 1666464484
transform 0 -1 16283 1 0 7672
box -88 -44 208 572
use nmos_5p043105899832103_64x8m81  nmos_5p043105899832103_64x8m81_1
timestamp 1666464484
transform 0 -1 11913 1 0 7672
box -88 -44 208 572
use pmos_1p2$$204216364_R90_64x8m81  pmos_1p2$$204216364_R90_64x8m81_0
timestamp 1666464484
transform 0 -1 20950 1 0 7703
box -296 -137 586 2646
use pmos_1p2$$204216364_R90_64x8m81  pmos_1p2$$204216364_R90_64x8m81_1
timestamp 1666464484
transform 0 -1 9245 1 0 7703
box -296 -137 586 2646
use pmos_1p2$$204217388_R90_64x8m81  pmos_1p2$$204217388_R90_64x8m81_0
timestamp 1666464484
transform 0 -1 11004 1 0 7703
box -295 -137 355 1454
use pmos_5p043105899832101_64x8m81  pmos_5p043105899832101_64x8m81_0
timestamp 1666464484
transform 0 -1 15304 1 0 7672
box -208 -120 328 1438
use pmos_5p043105899832101_64x8m81  pmos_5p043105899832101_64x8m81_1
timestamp 1666464484
transform 0 -1 17974 1 0 7672
box -208 -120 328 1438
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 2203 -1 0 7350
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_1
timestamp 1666464484
transform 0 -1 2203 -1 0 5550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_2
timestamp 1666464484
transform 0 -1 2203 -1 0 3750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_3
timestamp 1666464484
transform 0 -1 2203 -1 0 1950
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_4
timestamp 1666464484
transform 0 1 25566 -1 0 7350
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_5
timestamp 1666464484
transform 0 1 25566 -1 0 5550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_6
timestamp 1666464484
transform 0 1 25566 -1 0 3750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_64x8m81  pmoscap_W2_5_477_R270_64x8m81_7
timestamp 1666464484
transform 0 1 25566 -1 0 1950
box -60 -407 2159 5567
use pmoscap_W2_5_R270_64x8m81  pmoscap_W2_5_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 2203 -1 0 8250
box -60 -407 1259 3251
use pmoscap_W2_5_R270_64x8m81  pmoscap_W2_5_R270_64x8m81_1
timestamp 1666464484
transform 0 1 25566 -1 0 8250
box -60 -407 1259 3251
use xdec8_64x8m81  xdec8_64x8m81_0
timestamp 1666464484
transform 1 0 1726 0 1 0
box 0 -228 24219 7428
<< labels >>
rlabel metal3 s 27705 7640 27705 7640 4 DRWL
port 1 nsew
rlabel metal3 s 27705 5860 27705 5860 4 RWL[6]
port 2 nsew
rlabel metal3 s 27705 4060 27705 4060 4 RWL[4]
port 3 nsew
rlabel metal3 s 27705 2260 27705 2260 4 RWL[2]
port 4 nsew
rlabel metal3 s 27705 460 27705 460 4 RWL[0]
port 5 nsew
rlabel metal3 s 27705 1340 27705 1340 4 RWL[1]
port 6 nsew
rlabel metal3 s 27705 3140 27705 3140 4 RWL[3]
port 7 nsew
rlabel metal3 s 27705 4940 27705 4940 4 RWL[5]
port 8 nsew
rlabel metal3 s 27705 6740 27705 6740 4 RWL[7]
port 9 nsew
rlabel metal3 s 2556 5840 2556 5840 4 LWL[6]
port 10 nsew
rlabel metal3 s 2556 6760 2556 6760 4 LWL[7]
port 11 nsew
rlabel metal3 s 2556 1360 2556 1360 4 LWL[1]
port 12 nsew
rlabel metal3 s 2556 2240 2556 2240 4 LWL[2]
port 13 nsew
rlabel metal3 s 2556 3160 2556 3160 4 LWL[3]
port 14 nsew
rlabel metal3 s 2556 4040 2556 4040 4 LWL[4]
port 15 nsew
rlabel metal3 s 2556 4960 2556 4960 4 LWL[5]
port 16 nsew
rlabel metal3 s 64 4940 64 4940 4 LWL[5]
port 16 nsew
rlabel metal3 s 64 4060 64 4060 4 LWL[4]
port 15 nsew
rlabel metal3 s 64 3140 64 3140 4 LWL[3]
port 14 nsew
rlabel metal3 s 64 2260 64 2260 4 LWL[2]
port 13 nsew
rlabel metal3 s 64 1340 64 1340 4 LWL[1]
port 12 nsew
rlabel metal3 s 64 460 64 460 4 LWL[0]
port 17 nsew
rlabel metal3 s 64 5860 64 5860 4 LWL[6]
port 10 nsew
rlabel metal3 s 64 6740 64 6740 4 LWL[7]
port 11 nsew
rlabel metal3 s 2556 440 2556 440 4 LWL[0]
port 17 nsew
rlabel metal3 s 134 8100 134 8100 4 vss
port 18 nsew
rlabel metal3 s 134 7200 134 7200 4 vdd
port 19 nsew
rlabel metal3 s 64 7640 64 7640 4 DLWL
port 20 nsew
rlabel metal3 s 25149 6760 25149 6760 4 RWL[7]
port 9 nsew
rlabel metal3 s 25149 4960 25149 4960 4 RWL[5]
port 8 nsew
rlabel metal3 s 25149 3160 25149 3160 4 RWL[3]
port 7 nsew
rlabel metal3 s 25149 1360 25149 1360 4 RWL[1]
port 6 nsew
rlabel metal3 s 25149 440 25149 440 4 RWL[0]
port 5 nsew
rlabel metal3 s 25149 2240 25149 2240 4 RWL[2]
port 4 nsew
rlabel metal3 s 25149 4040 25149 4040 4 RWL[4]
port 3 nsew
rlabel metal3 s 25149 5840 25149 5840 4 RWL[6]
port 2 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 21 nsew
rlabel metal2 s 16947 -97 16947 -97 4 xa[7]
port 22 nsew
rlabel metal2 s 17324 -97 17324 -97 4 xa[6]
port 23 nsew
rlabel metal2 s 17702 -97 17702 -97 4 xa[5]
port 24 nsew
rlabel metal2 s 18080 -97 18080 -97 4 xa[4]
port 25 nsew
rlabel metal2 s 19591 -97 19591 -97 4 xa[0]
port 26 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 21 nsew
rlabel metal2 s 18457 -97 18457 -97 4 xa[3]
port 27 nsew
rlabel metal2 s 18835 -97 18835 -97 4 xa[2]
port 28 nsew
rlabel metal2 s 19213 -97 19213 -97 4 xa[1]
port 29 nsew
<< properties >>
string GDS_END 1864754
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1849354
<< end >>
