magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -30 363 88 436
rect 193 363 312 431
rect -30 -74 88 -1
rect 194 -74 312 -1
use nmos_5p04310589983263_64x8m81  nmos_5p04310589983263_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 432 408
<< properties >>
string GDS_END 9854
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 9476
<< end >>
