magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -19 248 19 253
rect -19 -248 -14 248
rect 14 -248 19 248
rect -19 -253 19 -248
<< via2 >>
rect -14 -248 14 248
<< metal3 >>
rect -19 248 19 253
rect -19 -248 -14 248
rect 14 -248 19 248
rect -19 -253 19 -248
<< properties >>
string GDS_END 569106
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 568334
<< end >>
