magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1878 1094
<< pwell >>
rect -86 -86 1878 453
<< mvnmos >>
rect 124 69 324 333
rect 572 69 772 333
rect 1020 69 1220 333
rect 1468 69 1668 333
<< mvpmos >>
rect 124 573 324 939
rect 572 573 772 939
rect 1020 573 1220 939
rect 1468 573 1668 939
<< mvndiff >>
rect 36 287 124 333
rect 36 147 49 287
rect 95 147 124 287
rect 36 69 124 147
rect 324 287 412 333
rect 324 147 353 287
rect 399 147 412 287
rect 324 69 412 147
rect 484 287 572 333
rect 484 147 497 287
rect 543 147 572 287
rect 484 69 572 147
rect 772 287 860 333
rect 772 147 801 287
rect 847 147 860 287
rect 772 69 860 147
rect 932 287 1020 333
rect 932 147 945 287
rect 991 147 1020 287
rect 932 69 1020 147
rect 1220 287 1308 333
rect 1220 147 1249 287
rect 1295 147 1308 287
rect 1220 69 1308 147
rect 1380 287 1468 333
rect 1380 147 1393 287
rect 1439 147 1468 287
rect 1380 69 1468 147
rect 1668 287 1756 333
rect 1668 147 1697 287
rect 1743 147 1756 287
rect 1668 69 1756 147
<< mvpdiff >>
rect 36 861 124 939
rect 36 721 49 861
rect 95 721 124 861
rect 36 573 124 721
rect 324 861 412 939
rect 324 721 353 861
rect 399 721 412 861
rect 324 573 412 721
rect 484 861 572 939
rect 484 721 497 861
rect 543 721 572 861
rect 484 573 572 721
rect 772 861 860 939
rect 772 721 801 861
rect 847 721 860 861
rect 772 573 860 721
rect 932 861 1020 939
rect 932 721 945 861
rect 991 721 1020 861
rect 932 573 1020 721
rect 1220 861 1308 939
rect 1220 721 1249 861
rect 1295 721 1308 861
rect 1220 573 1308 721
rect 1380 861 1468 939
rect 1380 721 1393 861
rect 1439 721 1468 861
rect 1380 573 1468 721
rect 1668 861 1756 939
rect 1668 721 1697 861
rect 1743 721 1756 861
rect 1668 573 1756 721
<< mvndiffc >>
rect 49 147 95 287
rect 353 147 399 287
rect 497 147 543 287
rect 801 147 847 287
rect 945 147 991 287
rect 1249 147 1295 287
rect 1393 147 1439 287
rect 1697 147 1743 287
<< mvpdiffc >>
rect 49 721 95 861
rect 353 721 399 861
rect 497 721 543 861
rect 801 721 847 861
rect 945 721 991 861
rect 1249 721 1295 861
rect 1393 721 1439 861
rect 1697 721 1743 861
<< polysilicon >>
rect 124 939 324 983
rect 572 939 772 983
rect 1020 939 1220 983
rect 1468 939 1668 983
rect 124 540 324 573
rect 124 494 265 540
rect 311 494 324 540
rect 124 481 324 494
rect 572 540 772 573
rect 572 494 713 540
rect 759 494 772 540
rect 572 481 772 494
rect 1020 540 1220 573
rect 1020 494 1161 540
rect 1207 494 1220 540
rect 1020 481 1220 494
rect 1468 540 1668 573
rect 1468 494 1609 540
rect 1655 494 1668 540
rect 1468 481 1668 494
rect 124 412 324 425
rect 124 366 137 412
rect 183 366 324 412
rect 124 333 324 366
rect 572 412 772 425
rect 572 366 585 412
rect 631 366 772 412
rect 572 333 772 366
rect 1020 412 1220 425
rect 1020 366 1033 412
rect 1079 366 1220 412
rect 1020 333 1220 366
rect 1468 412 1668 425
rect 1468 366 1481 412
rect 1527 366 1668 412
rect 1468 333 1668 366
rect 124 25 324 69
rect 572 25 772 69
rect 1020 25 1220 69
rect 1468 25 1668 69
<< polycontact >>
rect 265 494 311 540
rect 713 494 759 540
rect 1161 494 1207 540
rect 1609 494 1655 540
rect 137 366 183 412
rect 585 366 631 412
rect 1033 366 1079 412
rect 1481 366 1527 412
<< metal1 >>
rect 0 918 1792 1098
rect 49 861 95 872
rect 49 412 95 721
rect 353 861 399 918
rect 353 710 399 721
rect 497 861 543 872
rect 254 494 265 540
rect 311 494 399 540
rect 49 366 137 412
rect 183 366 194 412
rect 49 287 95 298
rect 49 90 95 147
rect 353 287 399 494
rect 497 412 543 721
rect 801 861 847 918
rect 801 710 847 721
rect 945 861 991 872
rect 702 494 713 540
rect 759 494 847 540
rect 497 366 585 412
rect 631 366 642 412
rect 353 136 399 147
rect 497 287 543 298
rect 497 90 543 147
rect 801 287 847 494
rect 945 412 991 721
rect 1249 861 1295 918
rect 1249 710 1295 721
rect 1393 861 1439 872
rect 1150 494 1161 540
rect 1207 494 1295 540
rect 945 366 1033 412
rect 1079 366 1090 412
rect 801 136 847 147
rect 945 287 991 298
rect 945 90 991 147
rect 1249 287 1295 494
rect 1393 412 1439 721
rect 1697 861 1743 918
rect 1697 710 1743 721
rect 1598 494 1609 540
rect 1655 494 1743 540
rect 1393 366 1481 412
rect 1527 366 1538 412
rect 1249 136 1295 147
rect 1393 287 1439 298
rect 1393 90 1439 147
rect 1697 287 1743 494
rect 1697 136 1743 147
rect 0 -90 1792 90
<< labels >>
flabel metal1 s 0 918 1792 1098 0 FreeSans 200 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 1393 90 1439 298 0 FreeSans 200 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 1697 710 1743 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 710 1295 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 710 847 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 710 399 918 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 945 90 991 298 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 298 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 298 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1792 90 1 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 1008
string GDS_END 769672
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 764158
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
