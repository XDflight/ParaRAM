magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 2128 844
rect 59 506 105 724
rect 273 552 319 675
rect 466 604 534 724
rect 594 632 1270 678
rect 594 552 640 632
rect 1320 586 1848 652
rect 273 506 640 552
rect 694 584 1848 586
rect 694 539 1370 584
rect 56 354 426 430
rect 472 244 536 506
rect 694 424 760 539
rect 1451 493 1670 538
rect 892 447 1670 493
rect 892 430 998 447
rect 594 354 760 424
rect 806 354 998 430
rect 1084 336 1395 397
rect 1534 382 1670 447
rect 1802 382 1848 584
rect 1898 506 1966 724
rect 1924 336 1996 456
rect 1084 333 1996 336
rect 1349 290 1996 333
rect 472 198 1720 244
rect 1794 242 1996 290
rect 262 60 330 127
rect 0 -60 2128 60
<< obsm1 >>
rect 36 173 426 219
rect 380 152 426 173
rect 380 106 1988 152
<< labels >>
rlabel metal1 s 1924 397 1996 456 6 A1
port 1 nsew default input
rlabel metal1 s 1924 336 1996 397 6 A1
port 1 nsew default input
rlabel metal1 s 1084 336 1395 397 6 A1
port 1 nsew default input
rlabel metal1 s 1084 333 1996 336 6 A1
port 1 nsew default input
rlabel metal1 s 1349 290 1996 333 6 A1
port 1 nsew default input
rlabel metal1 s 1794 242 1996 290 6 A1
port 1 nsew default input
rlabel metal1 s 1451 493 1670 538 6 A2
port 2 nsew default input
rlabel metal1 s 892 447 1670 493 6 A2
port 2 nsew default input
rlabel metal1 s 1534 430 1670 447 6 A2
port 2 nsew default input
rlabel metal1 s 892 430 998 447 6 A2
port 2 nsew default input
rlabel metal1 s 1534 382 1670 430 6 A2
port 2 nsew default input
rlabel metal1 s 806 382 998 430 6 A2
port 2 nsew default input
rlabel metal1 s 806 354 998 382 6 A2
port 2 nsew default input
rlabel metal1 s 1320 586 1848 652 6 A3
port 3 nsew default input
rlabel metal1 s 694 584 1848 586 6 A3
port 3 nsew default input
rlabel metal1 s 1802 539 1848 584 6 A3
port 3 nsew default input
rlabel metal1 s 694 539 1370 584 6 A3
port 3 nsew default input
rlabel metal1 s 1802 424 1848 539 6 A3
port 3 nsew default input
rlabel metal1 s 694 424 760 539 6 A3
port 3 nsew default input
rlabel metal1 s 1802 382 1848 424 6 A3
port 3 nsew default input
rlabel metal1 s 594 382 760 424 6 A3
port 3 nsew default input
rlabel metal1 s 594 354 760 382 6 A3
port 3 nsew default input
rlabel metal1 s 56 354 426 430 6 B
port 4 nsew default input
rlabel metal1 s 594 675 1270 678 6 ZN
port 5 nsew default output
rlabel metal1 s 594 632 1270 675 6 ZN
port 5 nsew default output
rlabel metal1 s 273 632 319 675 6 ZN
port 5 nsew default output
rlabel metal1 s 594 552 640 632 6 ZN
port 5 nsew default output
rlabel metal1 s 273 552 319 632 6 ZN
port 5 nsew default output
rlabel metal1 s 273 506 640 552 6 ZN
port 5 nsew default output
rlabel metal1 s 472 244 536 506 6 ZN
port 5 nsew default output
rlabel metal1 s 472 198 1720 244 6 ZN
port 5 nsew default output
rlabel metal1 s 0 724 2128 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1898 604 1966 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 466 604 534 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 604 105 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1898 506 1966 604 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 506 105 604 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 60 330 127 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2128 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2128 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 43126
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 38456
<< end >>
