magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 603 88 677
rect -31 -74 88 -1
use nmos_5p04310590878190_256x8m81  nmos_5p04310590878190_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 208 648
<< properties >>
string GDS_END 1063598
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1063348
<< end >>
