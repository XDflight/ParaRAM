magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 2998 870
rect -86 352 1922 377
rect 2678 352 2998 377
<< pwell >>
rect 1922 352 2678 377
rect -86 -86 2998 352
<< mvnmos >>
rect 124 68 244 232
rect 328 68 448 232
rect 552 68 672 232
rect 756 68 876 232
rect 980 68 1100 232
rect 1184 68 1304 232
rect 1408 68 1528 232
rect 1612 68 1732 232
rect 1816 68 1936 232
rect 2128 68 2248 232
rect 2352 68 2472 232
rect 2664 68 2784 232
<< mvpmos >>
rect 124 519 224 716
rect 328 519 428 716
rect 552 519 652 716
rect 756 519 856 716
rect 980 519 1080 716
rect 1184 519 1284 716
rect 1408 519 1508 716
rect 1612 519 1712 716
rect 1816 519 1916 716
rect 2128 519 2228 716
rect 2352 519 2452 716
rect 2664 519 2764 716
<< mvndiff >>
rect 1996 244 2068 257
rect 1996 232 2009 244
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 68 328 232
rect 448 127 552 232
rect 448 81 477 127
rect 523 81 552 127
rect 448 68 552 81
rect 672 68 756 232
rect 876 152 980 232
rect 876 106 905 152
rect 951 106 980 152
rect 876 68 980 106
rect 1100 68 1184 232
rect 1304 127 1408 232
rect 1304 81 1333 127
rect 1379 81 1408 127
rect 1304 68 1408 81
rect 1528 68 1612 232
rect 1732 68 1816 232
rect 1936 198 2009 232
rect 2055 232 2068 244
rect 2532 244 2604 257
rect 2532 232 2545 244
rect 2055 198 2128 232
rect 1936 68 2128 198
rect 2248 152 2352 232
rect 2248 106 2277 152
rect 2323 106 2352 152
rect 2248 68 2352 106
rect 2472 198 2545 232
rect 2591 232 2604 244
rect 2591 198 2664 232
rect 2472 68 2664 198
rect 2784 152 2872 232
rect 2784 106 2813 152
rect 2859 106 2872 152
rect 2784 68 2872 106
<< mvpdiff >>
rect 36 703 124 716
rect 36 563 49 703
rect 95 563 124 703
rect 36 519 124 563
rect 224 672 328 716
rect 224 532 253 672
rect 299 532 328 672
rect 224 519 328 532
rect 428 654 552 716
rect 428 608 457 654
rect 503 608 552 654
rect 428 519 552 608
rect 652 672 756 716
rect 652 532 681 672
rect 727 532 756 672
rect 652 519 756 532
rect 856 654 980 716
rect 856 608 885 654
rect 931 608 980 654
rect 856 519 980 608
rect 1080 672 1184 716
rect 1080 532 1109 672
rect 1155 532 1184 672
rect 1080 519 1184 532
rect 1284 654 1408 716
rect 1284 608 1313 654
rect 1359 608 1408 654
rect 1284 519 1408 608
rect 1508 672 1612 716
rect 1508 532 1537 672
rect 1583 532 1612 672
rect 1508 519 1612 532
rect 1712 654 1816 716
rect 1712 608 1741 654
rect 1787 608 1816 654
rect 1712 519 1816 608
rect 1916 672 2128 716
rect 1916 532 2009 672
rect 2055 532 2128 672
rect 1916 519 2128 532
rect 2228 654 2352 716
rect 2228 608 2257 654
rect 2303 608 2352 654
rect 2228 519 2352 608
rect 2452 672 2664 716
rect 2452 532 2545 672
rect 2591 532 2664 672
rect 2452 519 2664 532
rect 2764 703 2852 716
rect 2764 563 2793 703
rect 2839 563 2852 703
rect 2764 519 2852 563
<< mvndiffc >>
rect 49 173 95 219
rect 477 81 523 127
rect 905 106 951 152
rect 1333 81 1379 127
rect 2009 198 2055 244
rect 2277 106 2323 152
rect 2545 198 2591 244
rect 2813 106 2859 152
<< mvpdiffc >>
rect 49 563 95 703
rect 253 532 299 672
rect 457 608 503 654
rect 681 532 727 672
rect 885 608 931 654
rect 1109 532 1155 672
rect 1313 608 1359 654
rect 1537 532 1583 672
rect 1741 608 1787 654
rect 2009 532 2055 672
rect 2257 608 2303 654
rect 2545 532 2591 672
rect 2793 563 2839 703
<< polysilicon >>
rect 124 716 224 760
rect 328 716 428 760
rect 552 716 652 760
rect 756 716 856 760
rect 980 716 1080 760
rect 1184 716 1284 760
rect 1408 716 1508 760
rect 1612 716 1712 760
rect 1816 716 1916 760
rect 2128 716 2228 760
rect 2352 716 2452 760
rect 2664 716 2764 760
rect 124 415 224 519
rect 124 369 152 415
rect 198 369 224 415
rect 124 288 224 369
rect 328 394 428 519
rect 552 394 652 519
rect 328 348 652 394
rect 328 312 448 348
rect 124 232 244 288
rect 328 266 368 312
rect 414 266 448 312
rect 328 232 448 266
rect 552 312 652 348
rect 552 266 582 312
rect 628 288 652 312
rect 756 415 856 519
rect 756 369 789 415
rect 835 394 856 415
rect 980 415 1080 519
rect 980 394 1007 415
rect 835 369 1007 394
rect 1053 369 1080 415
rect 756 348 1080 369
rect 628 266 672 288
rect 552 232 672 266
rect 756 232 876 348
rect 980 288 1080 348
rect 1184 394 1284 519
rect 1408 394 1508 519
rect 1184 348 1508 394
rect 1184 312 1304 348
rect 980 232 1100 288
rect 1184 266 1222 312
rect 1268 266 1304 312
rect 1184 232 1304 266
rect 1408 312 1508 348
rect 1408 266 1441 312
rect 1487 288 1508 312
rect 1612 415 1712 519
rect 1612 369 1640 415
rect 1686 369 1712 415
rect 1612 288 1712 369
rect 1816 428 1916 519
rect 2128 428 2228 519
rect 2352 428 2452 519
rect 2664 428 2764 519
rect 1816 415 2764 428
rect 1816 369 1830 415
rect 2534 369 2764 415
rect 1816 356 2764 369
rect 1487 266 1528 288
rect 1408 232 1528 266
rect 1612 232 1732 288
rect 1816 232 1936 356
rect 2128 232 2248 356
rect 2352 232 2472 356
rect 2664 288 2764 356
rect 2664 232 2784 288
rect 124 24 244 68
rect 328 24 448 68
rect 552 24 672 68
rect 756 24 876 68
rect 980 24 1100 68
rect 1184 24 1304 68
rect 1408 24 1528 68
rect 1612 24 1732 68
rect 1816 24 1936 68
rect 2128 24 2248 68
rect 2352 24 2472 68
rect 2664 24 2784 68
<< polycontact >>
rect 152 369 198 415
rect 368 266 414 312
rect 582 266 628 312
rect 789 369 835 415
rect 1007 369 1053 415
rect 1222 266 1268 312
rect 1441 266 1487 312
rect 1640 369 1686 415
rect 1830 369 2534 415
<< metal1 >>
rect 0 724 2912 844
rect 49 703 95 724
rect 49 552 95 563
rect 242 532 253 672
rect 299 551 310 672
rect 457 654 503 724
rect 457 597 503 608
rect 670 551 681 672
rect 299 532 681 551
rect 727 551 738 672
rect 885 654 931 724
rect 885 597 931 608
rect 1098 551 1109 672
rect 727 532 1109 551
rect 1155 551 1166 672
rect 1313 654 1359 724
rect 1313 597 1359 608
rect 1526 551 1537 672
rect 1155 532 1537 551
rect 1583 551 1594 672
rect 1741 654 1787 724
rect 1741 597 1787 608
rect 1998 551 2009 672
rect 1583 532 2009 551
rect 2055 551 2066 672
rect 2257 654 2303 724
rect 2793 703 2839 724
rect 2257 597 2303 608
rect 2532 551 2545 672
rect 2055 532 2545 551
rect 2591 532 2670 672
rect 2793 552 2839 563
rect 242 476 2670 532
rect 130 415 1706 430
rect 130 369 152 415
rect 198 369 789 415
rect 835 369 1007 415
rect 1053 369 1640 415
rect 1686 369 1706 415
rect 130 358 1706 369
rect 1810 415 2534 426
rect 1810 369 1830 415
rect 1810 358 2534 369
rect 342 266 368 312
rect 414 266 582 312
rect 628 266 1222 312
rect 1268 266 1441 312
rect 1487 266 1508 312
rect 690 242 1132 266
rect 2594 244 2670 476
rect 36 173 49 219
rect 95 173 635 219
rect 589 152 635 173
rect 1227 173 1596 220
rect 1936 198 2009 244
rect 2055 198 2545 244
rect 2591 198 2670 244
rect 1227 152 1273 173
rect 464 81 477 127
rect 523 81 536 127
rect 589 106 905 152
rect 951 106 1273 152
rect 1550 152 1596 173
rect 464 60 536 81
rect 1320 81 1333 127
rect 1379 81 1392 127
rect 1550 106 2277 152
rect 2323 106 2813 152
rect 2859 106 2872 152
rect 1320 60 1392 81
rect 0 -60 2912 60
<< labels >>
flabel metal1 s 342 266 1508 312 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 2912 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1320 60 1392 127 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2532 551 2670 672 0 FreeSans 400 0 0 0 ZN
port 4 nsew default output
flabel metal1 s 1810 358 2534 426 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 130 358 1706 430 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 690 242 1132 266 1 A3
port 3 nsew default input
rlabel metal1 s 1998 551 2066 672 1 ZN
port 4 nsew default output
rlabel metal1 s 1526 551 1594 672 1 ZN
port 4 nsew default output
rlabel metal1 s 1098 551 1166 672 1 ZN
port 4 nsew default output
rlabel metal1 s 670 551 738 672 1 ZN
port 4 nsew default output
rlabel metal1 s 242 551 310 672 1 ZN
port 4 nsew default output
rlabel metal1 s 242 476 2670 551 1 ZN
port 4 nsew default output
rlabel metal1 s 2594 244 2670 476 1 ZN
port 4 nsew default output
rlabel metal1 s 1936 198 2670 244 1 ZN
port 4 nsew default output
rlabel metal1 s 2793 597 2839 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2257 597 2303 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1741 597 1787 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1313 597 1359 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 885 597 931 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 457 597 503 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 597 95 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2793 552 2839 597 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 552 95 597 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 464 60 536 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2912 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2912 784
string GDS_END 708848
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 702576
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
