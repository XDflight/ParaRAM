magic
tech gf180mcuC
magscale 1 5
timestamp 1667403444
<< checkpaint >>
rect 9200 9200 36500 36500
<< metal4 >>
rect 10200 24365 11700 35500
tri 11700 24365 12322 24987 sw
tri 10200 22932 11633 24365 ne
rect 11633 22932 12322 24365
tri 12322 22932 13755 24365 sw
tri 11633 20810 13755 22932 ne
tri 13755 20810 15877 22932 sw
tri 13755 18688 15877 20810 ne
tri 15877 18688 17999 20810 sw
tri 15877 16566 17999 18688 ne
tri 17999 16566 20121 18688 sw
tri 17999 14444 20121 16566 ne
tri 20121 14444 22243 16566 sw
tri 20121 12322 22243 14444 ne
tri 22243 12322 24365 14444 sw
tri 22243 10200 24365 12322 ne
tri 24365 11700 24987 12322 sw
rect 24365 10200 35500 11700
<< end >>
