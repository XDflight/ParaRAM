magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 2886 870
<< pwell >>
rect -86 -86 2886 352
<< mvnmos >>
rect 174 68 294 140
rect 398 68 518 140
rect 566 68 686 140
rect 1022 68 1142 140
rect 1190 68 1310 140
rect 1414 68 1534 140
rect 1582 68 1702 140
rect 2058 68 2178 141
rect 2226 68 2346 141
rect 2556 68 2676 232
<< mvpmos >>
rect 174 644 274 716
rect 398 644 498 716
rect 566 644 666 716
rect 1002 644 1102 716
rect 1170 644 1270 716
rect 1454 644 1554 716
rect 1622 644 1722 716
rect 2058 622 2158 694
rect 2226 622 2326 694
rect 2556 472 2656 716
<< mvndiff >>
rect 42 180 114 193
rect 42 134 55 180
rect 101 140 114 180
rect 746 200 818 213
rect 746 154 759 200
rect 805 154 818 200
rect 746 140 818 154
rect 101 134 174 140
rect 42 68 174 134
rect 294 127 398 140
rect 294 81 323 127
rect 369 81 398 127
rect 294 68 398 81
rect 518 68 566 140
rect 686 68 818 140
rect 890 200 962 213
rect 890 154 903 200
rect 949 154 962 200
rect 890 140 962 154
rect 1762 200 1834 213
rect 1762 154 1775 200
rect 1821 154 1834 200
rect 1762 140 1834 154
rect 890 68 1022 140
rect 1142 68 1190 140
rect 1310 127 1414 140
rect 1310 81 1339 127
rect 1385 81 1414 127
rect 1310 68 1414 81
rect 1534 68 1582 140
rect 1702 68 1834 140
rect 1926 200 1998 213
rect 1926 154 1939 200
rect 1985 154 1998 200
rect 1926 141 1998 154
rect 2476 141 2556 232
rect 1926 68 2058 141
rect 2178 68 2226 141
rect 2346 127 2556 141
rect 2346 81 2423 127
rect 2469 81 2556 127
rect 2346 68 2556 81
rect 2676 192 2764 232
rect 2676 146 2705 192
rect 2751 146 2764 192
rect 2676 68 2764 146
<< mvpdiff >>
rect 42 644 174 716
rect 274 703 398 716
rect 274 657 303 703
rect 349 657 398 703
rect 274 644 398 657
rect 498 644 566 716
rect 666 644 798 716
rect 42 621 114 644
rect 42 575 55 621
rect 101 575 114 621
rect 42 562 114 575
rect 726 621 798 644
rect 726 575 739 621
rect 785 575 798 621
rect 726 562 798 575
rect 870 644 1002 716
rect 1102 644 1170 716
rect 1270 703 1454 716
rect 1270 657 1299 703
rect 1345 657 1454 703
rect 1270 644 1454 657
rect 1554 644 1622 716
rect 1722 644 1854 716
rect 2476 694 2556 716
rect 870 621 942 644
rect 870 575 883 621
rect 929 575 942 621
rect 870 562 942 575
rect 1782 621 1854 644
rect 1782 575 1795 621
rect 1841 575 1854 621
rect 1782 562 1854 575
rect 1926 622 2058 694
rect 2158 622 2226 694
rect 2326 681 2556 694
rect 2326 635 2355 681
rect 2401 635 2556 681
rect 2326 622 2556 635
rect 1926 621 1998 622
rect 1926 575 1939 621
rect 1985 575 1998 621
rect 1926 562 1998 575
rect 2476 472 2556 622
rect 2656 639 2744 716
rect 2656 593 2685 639
rect 2731 593 2744 639
rect 2656 531 2744 593
rect 2656 485 2685 531
rect 2731 485 2744 531
rect 2656 472 2744 485
<< mvndiffc >>
rect 55 134 101 180
rect 759 154 805 200
rect 323 81 369 127
rect 903 154 949 200
rect 1775 154 1821 200
rect 1339 81 1385 127
rect 1939 154 1985 200
rect 2423 81 2469 127
rect 2705 146 2751 192
<< mvpdiffc >>
rect 303 657 349 703
rect 55 575 101 621
rect 739 575 785 621
rect 1299 657 1345 703
rect 883 575 929 621
rect 1795 575 1841 621
rect 2355 635 2401 681
rect 1939 575 1985 621
rect 2685 593 2731 639
rect 2685 485 2731 531
<< polysilicon >>
rect 174 716 274 760
rect 398 716 498 760
rect 566 716 666 760
rect 1002 716 1102 760
rect 1170 716 1270 760
rect 1454 716 1554 760
rect 1622 716 1722 760
rect 174 303 274 644
rect 174 257 187 303
rect 233 257 274 303
rect 174 184 274 257
rect 398 483 498 644
rect 566 483 666 644
rect 2058 694 2158 738
rect 2226 694 2326 738
rect 2556 716 2656 760
rect 398 470 666 483
rect 398 424 411 470
rect 457 424 591 470
rect 637 424 666 470
rect 398 411 666 424
rect 398 184 498 411
rect 566 184 666 411
rect 1002 371 1102 644
rect 1170 371 1270 644
rect 1002 350 1270 371
rect 1002 304 1015 350
rect 1061 304 1270 350
rect 1002 290 1270 304
rect 174 140 294 184
rect 398 140 518 184
rect 566 140 686 184
rect 1022 140 1142 290
rect 1190 184 1270 290
rect 1454 371 1554 644
rect 1622 371 1722 644
rect 1454 350 1722 371
rect 1454 304 1467 350
rect 1607 304 1722 350
rect 1454 290 1722 304
rect 2058 377 2158 622
rect 2226 377 2326 622
rect 2058 364 2326 377
rect 2058 318 2071 364
rect 2211 318 2326 364
rect 2058 305 2326 318
rect 1454 184 1534 290
rect 1190 140 1310 184
rect 1414 140 1534 184
rect 1582 140 1702 290
rect 2058 185 2158 305
rect 2226 185 2326 305
rect 2556 325 2656 472
rect 2556 279 2569 325
rect 2615 323 2656 325
rect 2615 279 2676 323
rect 2556 232 2676 279
rect 2058 141 2178 185
rect 2226 141 2346 185
rect 174 24 294 68
rect 398 24 518 68
rect 566 24 686 68
rect 1022 24 1142 68
rect 1190 24 1310 68
rect 1414 24 1534 68
rect 1582 24 1702 68
rect 2058 24 2178 68
rect 2226 24 2346 68
rect 2556 24 2676 68
<< polycontact >>
rect 187 257 233 303
rect 411 424 457 470
rect 591 424 637 470
rect 1015 304 1061 350
rect 1467 304 1607 350
rect 2071 318 2211 364
rect 2569 279 2615 325
<< metal1 >>
rect 0 724 2800 844
rect 292 703 360 724
rect 292 657 303 703
rect 349 657 360 703
rect 1288 703 1356 724
rect 1288 657 1299 703
rect 1345 657 1356 703
rect 2344 681 2412 724
rect 2344 635 2355 681
rect 2401 635 2412 681
rect 739 621 785 632
rect 1775 621 1852 632
rect 44 575 55 621
rect 101 575 112 621
rect 44 481 112 575
rect 872 575 883 621
rect 929 575 1153 621
rect 44 470 648 481
rect 44 424 411 470
rect 457 424 591 470
rect 637 424 648 470
rect 44 413 648 424
rect 44 180 112 413
rect 739 361 785 575
rect 739 350 1061 361
rect 181 303 666 320
rect 181 257 187 303
rect 233 257 666 303
rect 181 240 666 257
rect 739 304 1015 350
rect 739 293 1061 304
rect 1107 350 1153 575
rect 1775 575 1795 621
rect 1841 575 1852 621
rect 1775 393 1852 575
rect 1939 621 1985 632
rect 1939 493 1985 575
rect 2674 593 2685 639
rect 2731 593 2751 639
rect 2674 542 2751 593
rect 2393 531 2751 542
rect 1939 447 2333 493
rect 2393 485 2685 531
rect 2731 485 2751 531
rect 2393 466 2751 485
rect 1775 364 2211 393
rect 1107 304 1467 350
rect 1607 304 1618 350
rect 1775 318 2071 364
rect 1775 307 2211 318
rect 2269 325 2333 447
rect 44 134 55 180
rect 101 134 112 180
rect 739 200 816 293
rect 1107 200 1153 304
rect 739 154 759 200
rect 805 154 816 200
rect 892 154 903 200
rect 949 154 1153 200
rect 1775 200 1821 307
rect 2269 279 2569 325
rect 2615 279 2626 325
rect 2269 211 2333 279
rect 1775 143 1821 154
rect 1939 200 2333 211
rect 1985 154 2333 200
rect 1939 143 2333 154
rect 2705 192 2751 466
rect 2423 127 2469 138
rect 2705 135 2751 146
rect 312 81 323 127
rect 369 81 380 127
rect 312 60 380 81
rect 1328 81 1339 127
rect 1385 81 1396 127
rect 1328 60 1396 81
rect 2423 60 2469 81
rect 0 -60 2800 60
<< labels >>
flabel metal1 s 2674 542 2751 639 0 FreeSans 400 0 0 0 Z
port 2 nsew default output
flabel metal1 s 2423 127 2469 138 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 181 240 666 320 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 724 2800 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 2393 466 2751 542 1 Z
port 2 nsew default output
rlabel metal1 s 2705 135 2751 466 1 Z
port 2 nsew default output
rlabel metal1 s 2344 657 2412 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1288 657 1356 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 292 657 360 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2344 635 2412 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2423 60 2469 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1328 60 1396 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 312 60 380 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2800 60 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2800 784
string GDS_END 1088680
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1083428
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
