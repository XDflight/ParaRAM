magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 60123 842 60142
rect -42 -23 -23 60123
rect 823 -23 842 60123
rect -42 -42 842 -23
<< psubdiffcont >>
rect -23 -23 823 60123
<< metal1 >>
rect -34 60123 834 60134
rect -34 -23 -23 60123
rect 823 -23 834 60123
rect -34 -34 834 -23
<< properties >>
string GDS_END 1904704
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1557756
<< end >>
