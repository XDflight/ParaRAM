magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 2409
<< polysilicon >>
rect -31 2268 89 2330
rect -30 -74 88 0
use pmos_5p04310590548772_128x8m81  pmos_5p04310590548772_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 2388
<< properties >>
string GDS_END 344024
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 343710
<< end >>
