magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 792 595
<< polysilicon >>
rect -31 454 89 527
rect 193 454 313 527
rect 417 454 537 527
rect -31 -73 89 -1
rect 193 -73 313 -1
rect 417 -73 537 -1
use pmos_5p04310591302013_512x8m81  pmos_5p04310591302013_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 776 574
<< properties >>
string GDS_END 337020
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 336450
<< end >>
