magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 5126 1094
<< pwell >>
rect -86 -86 5126 453
<< mvnmos >>
rect 139 196 259 314
rect 363 196 483 314
rect 531 196 651 314
rect 755 196 875 314
rect 923 196 1043 314
rect 1323 164 1443 322
rect 1547 164 1667 322
rect 1915 174 2035 292
rect 2139 174 2259 292
rect 2307 174 2427 292
rect 2575 215 2695 333
rect 2759 215 2879 333
rect 2983 215 3103 333
rect 3207 215 3327 333
rect 3743 215 3863 333
rect 3927 215 4047 333
rect 4187 69 4307 333
rect 4572 69 4692 333
rect 4796 69 4916 333
<< mvpmos >>
rect 159 644 259 844
rect 383 644 483 844
rect 541 644 641 844
rect 755 644 855 844
rect 903 644 1003 844
rect 1343 573 1443 849
rect 1547 573 1647 849
rect 1925 582 2025 782
rect 2139 582 2239 782
rect 2327 582 2427 782
rect 2575 582 2675 782
rect 2779 582 2879 782
rect 3207 573 3307 773
rect 3415 573 3515 773
rect 3763 623 3863 823
rect 3967 623 4067 823
rect 4207 573 4307 939
rect 4592 573 4692 939
rect 4796 573 4896 939
<< mvndiff >>
rect 51 285 139 314
rect 51 239 64 285
rect 110 239 139 285
rect 51 196 139 239
rect 259 285 363 314
rect 259 239 288 285
rect 334 239 363 285
rect 259 196 363 239
rect 483 196 531 314
rect 651 285 755 314
rect 651 239 680 285
rect 726 239 755 285
rect 651 196 755 239
rect 875 196 923 314
rect 1043 196 1163 314
rect 1103 116 1163 196
rect 1235 309 1323 322
rect 1235 263 1248 309
rect 1294 263 1323 309
rect 1235 164 1323 263
rect 1443 223 1547 322
rect 1443 177 1472 223
rect 1518 177 1547 223
rect 1443 164 1547 177
rect 1667 285 1755 322
rect 2495 292 2575 333
rect 1667 239 1696 285
rect 1742 239 1755 285
rect 1667 164 1755 239
rect 1827 233 1915 292
rect 1827 187 1840 233
rect 1886 187 1915 233
rect 1827 174 1915 187
rect 2035 279 2139 292
rect 2035 233 2064 279
rect 2110 233 2139 279
rect 2035 174 2139 233
rect 2259 174 2307 292
rect 2427 233 2575 292
rect 2427 187 2456 233
rect 2502 215 2575 233
rect 2695 215 2759 333
rect 2879 285 2983 333
rect 2879 239 2908 285
rect 2954 239 2983 285
rect 2879 215 2983 239
rect 3103 285 3207 333
rect 3103 239 3132 285
rect 3178 239 3207 285
rect 3103 215 3207 239
rect 3327 320 3415 333
rect 3327 274 3356 320
rect 3402 274 3415 320
rect 3327 215 3415 274
rect 2502 187 2515 215
rect 2427 174 2515 187
rect 1096 114 1163 116
rect 1096 104 1168 114
rect 1096 58 1109 104
rect 1155 58 1168 104
rect 1096 45 1168 58
rect 3621 320 3743 333
rect 3621 274 3634 320
rect 3680 274 3743 320
rect 3621 215 3743 274
rect 3863 215 3927 333
rect 4047 285 4187 333
rect 4047 239 4076 285
rect 4122 239 4187 285
rect 4047 215 4187 239
rect 4107 69 4187 215
rect 4307 320 4395 333
rect 4307 180 4336 320
rect 4382 180 4395 320
rect 4307 69 4395 180
rect 4484 222 4572 333
rect 4484 82 4497 222
rect 4543 82 4572 222
rect 4484 69 4572 82
rect 4692 320 4796 333
rect 4692 180 4721 320
rect 4767 180 4796 320
rect 4692 69 4796 180
rect 4916 222 5004 333
rect 4916 82 4945 222
rect 4991 82 5004 222
rect 4916 69 5004 82
<< mvpdiff >>
rect 71 799 159 844
rect 71 659 84 799
rect 130 659 159 799
rect 71 644 159 659
rect 259 831 383 844
rect 259 691 288 831
rect 334 691 383 831
rect 259 644 383 691
rect 483 644 541 844
rect 641 831 755 844
rect 641 691 680 831
rect 726 691 755 831
rect 641 644 755 691
rect 855 644 903 844
rect 1003 809 1091 844
rect 1003 763 1032 809
rect 1078 763 1091 809
rect 1003 644 1091 763
rect 1255 632 1343 849
rect 1255 586 1268 632
rect 1314 586 1343 632
rect 1255 573 1343 586
rect 1443 829 1547 849
rect 1443 783 1472 829
rect 1518 783 1547 829
rect 1443 573 1547 783
rect 1647 726 1735 849
rect 4127 823 4207 939
rect 1647 586 1676 726
rect 1722 586 1735 726
rect 1647 573 1735 586
rect 1837 769 1925 782
rect 1837 629 1850 769
rect 1896 629 1925 769
rect 1837 582 1925 629
rect 2025 735 2139 782
rect 2025 595 2064 735
rect 2110 595 2139 735
rect 2025 582 2139 595
rect 2239 582 2327 782
rect 2427 769 2575 782
rect 2427 723 2456 769
rect 2502 723 2575 769
rect 2427 582 2575 723
rect 2675 735 2779 782
rect 2675 595 2704 735
rect 2750 595 2779 735
rect 2675 582 2779 595
rect 2879 769 2967 782
rect 3675 810 3763 823
rect 2879 723 2908 769
rect 2954 723 2967 769
rect 2879 582 2967 723
rect 3119 726 3207 773
rect 3119 586 3132 726
rect 3178 586 3207 726
rect 3119 573 3207 586
rect 3307 758 3415 773
rect 3307 618 3336 758
rect 3382 618 3415 758
rect 3307 573 3415 618
rect 3515 758 3603 773
rect 3515 618 3544 758
rect 3590 618 3603 758
rect 3675 670 3688 810
rect 3734 670 3763 810
rect 3675 623 3763 670
rect 3863 799 3967 823
rect 3863 659 3892 799
rect 3938 659 3967 799
rect 3863 623 3967 659
rect 4067 799 4207 823
rect 4067 659 4096 799
rect 4142 659 4207 799
rect 4067 623 4207 659
rect 3515 573 3603 618
rect 4127 573 4207 623
rect 4307 799 4395 939
rect 4307 659 4336 799
rect 4382 659 4395 799
rect 4307 573 4395 659
rect 4504 799 4592 939
rect 4504 659 4517 799
rect 4563 659 4592 799
rect 4504 573 4592 659
rect 4692 799 4796 939
rect 4692 659 4721 799
rect 4767 659 4796 799
rect 4692 573 4796 659
rect 4896 799 4984 939
rect 4896 659 4925 799
rect 4971 659 4984 799
rect 4896 573 4984 659
<< mvndiffc >>
rect 64 239 110 285
rect 288 239 334 285
rect 680 239 726 285
rect 1248 263 1294 309
rect 1472 177 1518 223
rect 1696 239 1742 285
rect 1840 187 1886 233
rect 2064 233 2110 279
rect 2456 187 2502 233
rect 2908 239 2954 285
rect 3132 239 3178 285
rect 3356 274 3402 320
rect 1109 58 1155 104
rect 3634 274 3680 320
rect 4076 239 4122 285
rect 4336 180 4382 320
rect 4497 82 4543 222
rect 4721 180 4767 320
rect 4945 82 4991 222
<< mvpdiffc >>
rect 84 659 130 799
rect 288 691 334 831
rect 680 691 726 831
rect 1032 763 1078 809
rect 1268 586 1314 632
rect 1472 783 1518 829
rect 1676 586 1722 726
rect 1850 629 1896 769
rect 2064 595 2110 735
rect 2456 723 2502 769
rect 2704 595 2750 735
rect 2908 723 2954 769
rect 3132 586 3178 726
rect 3336 618 3382 758
rect 3544 618 3590 758
rect 3688 670 3734 810
rect 3892 659 3938 799
rect 4096 659 4142 799
rect 4336 659 4382 799
rect 4517 659 4563 799
rect 4721 659 4767 799
rect 4925 659 4971 799
<< polysilicon >>
rect 159 936 1003 976
rect 159 844 259 936
rect 383 844 483 888
rect 541 844 641 888
rect 755 844 855 888
rect 903 844 1003 936
rect 1547 936 2239 976
rect 1343 849 1443 893
rect 1547 849 1647 936
rect 2139 861 2239 936
rect 159 510 259 644
rect 159 464 172 510
rect 218 464 259 510
rect 159 358 259 464
rect 383 510 483 644
rect 383 464 396 510
rect 442 464 483 510
rect 383 358 483 464
rect 541 510 641 644
rect 541 464 576 510
rect 622 464 641 510
rect 541 451 641 464
rect 755 510 855 644
rect 903 600 1003 644
rect 1925 782 2025 826
rect 2139 815 2180 861
rect 2226 815 2239 861
rect 2779 913 3863 953
rect 4207 939 4307 983
rect 4592 939 4692 983
rect 4796 939 4896 983
rect 2139 782 2239 815
rect 2327 782 2427 826
rect 2575 782 2675 826
rect 2779 782 2879 913
rect 3207 852 3307 865
rect 3207 806 3220 852
rect 3266 806 3307 852
rect 3763 823 3863 913
rect 3967 823 4067 867
rect 3207 773 3307 806
rect 3415 773 3515 817
rect 755 464 768 510
rect 814 464 855 510
rect 755 358 855 464
rect 923 510 1043 523
rect 923 464 936 510
rect 982 464 1043 510
rect 139 314 259 358
rect 363 314 483 358
rect 531 314 651 358
rect 755 314 875 358
rect 923 314 1043 464
rect 1343 510 1443 573
rect 1343 464 1384 510
rect 1430 464 1443 510
rect 1343 366 1443 464
rect 1323 322 1443 366
rect 1547 418 1647 573
rect 1925 510 2025 582
rect 2139 538 2239 582
rect 2327 549 2427 582
rect 1925 464 1938 510
rect 1984 490 2025 510
rect 2327 503 2368 549
rect 2414 503 2427 549
rect 1984 464 2259 490
rect 1925 418 2259 464
rect 1547 372 1560 418
rect 1606 372 1647 418
rect 1547 366 1647 372
rect 2139 371 2259 418
rect 1547 322 1667 366
rect 139 104 259 196
rect 363 152 483 196
rect 531 104 651 196
rect 755 152 875 196
rect 923 152 1043 196
rect 1915 292 2035 336
rect 2139 325 2180 371
rect 2226 325 2259 371
rect 2327 336 2427 503
rect 2139 292 2259 325
rect 2307 292 2427 336
rect 2575 457 2675 582
rect 2575 411 2588 457
rect 2634 411 2675 457
rect 2575 377 2675 411
rect 2779 377 2879 582
rect 3207 377 3307 573
rect 3415 529 3515 573
rect 2575 333 2695 377
rect 2759 333 2879 377
rect 2983 333 3103 377
rect 3207 333 3327 377
rect 1323 120 1443 164
rect 139 32 651 104
rect 1547 104 1667 164
rect 1915 104 2035 174
rect 2139 130 2259 174
rect 2307 130 2427 174
rect 2575 171 2695 215
rect 2759 171 2879 215
rect 2983 182 3103 215
rect 2983 136 2996 182
rect 3042 136 3103 182
rect 3207 171 3327 215
rect 1547 32 2035 104
rect 2983 123 3103 136
rect 3475 123 3515 529
rect 3763 510 3863 623
rect 3763 464 3776 510
rect 3822 464 3863 510
rect 3763 377 3863 464
rect 3967 510 4067 623
rect 3967 464 4008 510
rect 4054 464 4067 510
rect 3967 451 4067 464
rect 4207 510 4307 573
rect 4207 464 4220 510
rect 4266 464 4307 510
rect 3967 377 4047 451
rect 4207 377 4307 464
rect 4592 510 4692 573
rect 4592 464 4605 510
rect 4651 465 4692 510
rect 4796 465 4896 573
rect 4651 464 4896 465
rect 4592 393 4896 464
rect 4592 377 4692 393
rect 3743 333 3863 377
rect 3927 333 4047 377
rect 4187 333 4307 377
rect 4572 333 4692 377
rect 4796 377 4896 393
rect 4796 333 4916 377
rect 3743 171 3863 215
rect 3927 171 4047 215
rect 2983 51 3515 123
rect 4187 25 4307 69
rect 4572 25 4692 69
rect 4796 25 4916 69
<< polycontact >>
rect 172 464 218 510
rect 396 464 442 510
rect 576 464 622 510
rect 2180 815 2226 861
rect 3220 806 3266 852
rect 768 464 814 510
rect 936 464 982 510
rect 1384 464 1430 510
rect 1938 464 1984 510
rect 2368 503 2414 549
rect 1560 372 1606 418
rect 2180 325 2226 371
rect 2588 411 2634 457
rect 2996 136 3042 182
rect 3776 464 3822 510
rect 4008 464 4054 510
rect 4220 464 4266 510
rect 4605 464 4651 510
<< metal1 >>
rect 0 918 5040 1098
rect 288 831 334 918
rect 84 799 130 810
rect 288 680 334 691
rect 680 831 726 842
rect 1032 809 1078 918
rect 1472 829 1518 918
rect 2180 861 2226 872
rect 1472 772 1518 783
rect 1564 783 1896 829
rect 1032 752 1078 763
rect 1121 726 1444 735
rect 1564 726 1610 783
rect 1850 769 1896 783
rect 726 706 994 726
rect 1121 706 1610 726
rect 726 691 1610 706
rect 680 689 1610 691
rect 680 680 1164 689
rect 1416 680 1610 689
rect 1676 726 1722 737
rect 956 660 1164 680
rect 84 634 130 659
rect 1268 634 1314 643
rect 84 614 918 634
rect 1268 632 1630 634
rect 84 588 982 614
rect 142 510 306 542
rect 142 464 172 510
rect 218 464 306 510
rect 366 510 530 542
rect 366 464 396 510
rect 442 464 530 510
rect 576 510 622 588
rect 880 568 982 588
rect 1314 588 1630 632
rect 1268 575 1314 586
rect 576 418 622 464
rect 64 372 622 418
rect 702 510 814 542
rect 702 464 768 510
rect 64 285 110 372
rect 702 354 814 464
rect 936 510 982 568
rect 1373 510 1538 542
rect 1373 464 1384 510
rect 1430 464 1538 510
rect 936 453 982 464
rect 1584 418 1630 588
rect 1248 372 1560 418
rect 1606 372 1630 418
rect 1850 618 1896 629
rect 2064 735 2110 746
rect 1676 510 1722 586
rect 2180 666 2226 815
rect 2456 769 2502 918
rect 2456 712 2502 723
rect 2548 792 2862 838
rect 2548 666 2594 792
rect 2180 620 2594 666
rect 2704 735 2750 746
rect 1676 464 1938 510
rect 1984 464 1995 510
rect 1248 309 1294 372
rect 64 228 110 239
rect 288 285 334 296
rect 288 90 334 239
rect 680 285 726 296
rect 1248 252 1294 263
rect 1340 280 1610 326
rect 680 207 726 239
rect 680 206 1238 207
rect 1340 206 1386 280
rect 680 161 1386 206
rect 1228 160 1386 161
rect 1472 223 1518 234
rect 1109 104 1155 115
rect 0 58 1109 90
rect 1472 90 1518 177
rect 1564 182 1610 280
rect 1676 285 1742 464
rect 1676 239 1696 285
rect 2064 463 2110 595
rect 2816 666 2862 792
rect 2908 769 2954 918
rect 2908 712 2954 723
rect 3040 852 3266 863
rect 3040 806 3220 852
rect 3040 795 3266 806
rect 3688 810 3734 918
rect 3040 666 3086 795
rect 3336 758 3382 769
rect 2816 620 3086 666
rect 3132 726 3178 737
rect 2704 549 2750 595
rect 3132 549 3178 586
rect 2357 503 2368 549
rect 2414 503 3178 549
rect 2064 457 2334 463
rect 2064 417 2588 457
rect 2064 279 2110 417
rect 2311 411 2588 417
rect 2634 411 2645 457
rect 2169 325 2180 371
rect 2226 365 2237 371
rect 2226 325 2594 365
rect 2169 319 2594 325
rect 1676 228 1742 239
rect 1840 233 1886 244
rect 2064 222 2110 233
rect 2456 233 2502 244
rect 1840 182 1886 187
rect 1564 136 1886 182
rect 2456 90 2502 187
rect 2548 182 2594 319
rect 2908 285 2954 503
rect 3336 423 3382 618
rect 3544 758 3590 769
rect 3688 659 3734 670
rect 3892 799 3938 810
rect 3544 613 3590 618
rect 3892 613 3938 659
rect 4096 799 4142 918
rect 4096 648 4142 659
rect 4336 799 4382 810
rect 3544 567 3938 613
rect 4336 602 4382 659
rect 4517 799 4563 918
rect 4517 648 4563 659
rect 4721 799 4786 810
rect 4767 659 4786 799
rect 3264 377 3382 423
rect 3264 296 3310 377
rect 3634 331 3680 567
rect 4008 556 4651 602
rect 2908 228 2954 239
rect 3132 285 3310 296
rect 3178 239 3310 285
rect 3356 320 3680 331
rect 3402 274 3634 320
rect 3356 263 3680 274
rect 3726 510 3822 521
rect 3726 464 3776 510
rect 3726 453 3822 464
rect 4008 510 4054 556
rect 4008 453 4054 464
rect 4100 464 4220 510
rect 4266 464 4277 510
rect 3726 242 3778 453
rect 4100 388 4146 464
rect 3824 342 4146 388
rect 3132 228 3310 239
rect 3264 196 3310 228
rect 3824 196 3870 342
rect 4336 320 4382 556
rect 4605 510 4651 556
rect 4605 453 4651 464
rect 2548 136 2996 182
rect 3042 136 3053 182
rect 3264 150 3870 196
rect 4076 285 4122 296
rect 4076 90 4122 239
rect 4721 320 4786 659
rect 4925 799 4971 918
rect 4925 648 4971 659
rect 4336 169 4382 180
rect 4497 222 4543 233
rect 1155 82 4497 90
rect 4767 180 4786 320
rect 4721 169 4786 180
rect 4945 222 4991 233
rect 4543 82 4945 90
rect 4991 82 5040 90
rect 1155 58 5040 82
rect 0 -90 5040 58
<< labels >>
flabel metal1 s 1373 464 1538 542 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 702 354 814 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4721 169 4786 810 0 FreeSans 200 0 0 0 Q
port 6 nsew default output
flabel metal1 s 142 464 306 542 0 FreeSans 200 0 0 0 SE
port 2 nsew default input
flabel metal1 s 3726 453 3822 521 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 366 464 530 542 0 FreeSans 200 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 918 5040 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 4076 244 4122 296 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3726 242 3778 453 1 SETN
port 3 nsew default input
rlabel metal1 s 4925 772 4971 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 772 4563 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 772 4142 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3688 772 3734 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2908 772 2954 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2456 772 2502 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1472 772 1518 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1032 772 1078 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 288 772 334 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4925 752 4971 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 752 4563 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 752 4142 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3688 752 3734 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2908 752 2954 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2456 752 2502 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1032 752 1078 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 288 752 334 772 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4925 712 4971 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 712 4563 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 712 4142 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3688 712 3734 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2908 712 2954 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2456 712 2502 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 288 712 334 752 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4925 680 4971 712 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 680 4563 712 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 680 4142 712 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3688 680 3734 712 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 288 680 334 712 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4925 659 4971 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 659 4563 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 659 4142 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3688 659 3734 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4925 648 4971 659 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4517 648 4563 659 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4096 648 4142 659 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 288 244 334 296 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4076 234 4122 244 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2456 234 2502 244 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 288 234 334 244 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4076 233 4122 234 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2456 233 2502 234 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1472 233 1518 234 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 288 233 334 234 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4945 115 4991 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4497 115 4543 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4076 115 4122 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2456 115 2502 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1472 115 1518 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 288 115 334 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4945 90 4991 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4497 90 4543 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4076 90 4122 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2456 90 2502 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1472 90 1518 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1109 90 1155 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 288 90 334 115 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5040 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5040 1008
string GDS_END 420272
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 408510
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
