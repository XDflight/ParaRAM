magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 3406
<< polysilicon >>
rect -31 3265 88 3338
rect -31 -73 88 -1
use pmos_5p04310589983274_64x8m81  pmos_5p04310589983274_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 3386
<< properties >>
string GDS_END 153262
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 152948
<< end >>
