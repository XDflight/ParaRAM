magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -170 353 170 393
rect -170 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -170 135 170 301
rect -170 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -170 -83 170 83
rect -170 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -170 -301 170 -135
rect -170 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -170 -393 170 -353
<< via1 >>
rect -132 301 -80 353
rect 80 301 132 353
rect -132 83 -80 135
rect 80 83 132 135
rect -132 -135 -80 -83
rect 80 -135 132 -83
rect -132 -353 -80 -301
rect 80 -353 132 -301
<< metal2 >>
rect -169 353 170 393
rect -169 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -169 135 170 301
rect -169 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -169 -83 170 83
rect -169 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -169 -301 170 -135
rect -169 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -169 -393 170 -353
<< properties >>
string GDS_END 1115664
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1115020
<< end >>
