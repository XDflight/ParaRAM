magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 273 88 346
rect -31 -73 88 0
use nmos_5p04310591302040_512x8m81  nmos_5p04310591302040_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 208 318
<< properties >>
string GDS_END 218070
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 217820
<< end >>
