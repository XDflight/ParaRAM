magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 288
<< mvndiff >>
rect -88 275 0 288
rect -88 229 -75 275
rect -29 229 0 275
rect -88 167 0 229
rect -88 121 -75 167
rect -29 121 0 167
rect -88 59 0 121
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 275 208 288
rect 120 229 149 275
rect 195 229 208 275
rect 120 167 208 229
rect 120 121 149 167
rect 195 121 208 167
rect 120 59 208 121
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 229 -29 275
rect -75 121 -29 167
rect -75 13 -29 59
rect 149 229 195 275
rect 149 121 195 167
rect 149 13 195 59
<< polysilicon >>
rect 0 288 120 332
rect 0 -44 120 0
<< metal1 >>
rect -75 275 -29 288
rect -75 167 -29 229
rect -75 59 -29 121
rect -75 0 -29 13
rect 149 275 195 288
rect 149 167 195 229
rect 149 59 195 121
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 144 -52 144 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 144 172 144 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 273068
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 271788
<< end >>
