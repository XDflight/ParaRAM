magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -381 355 381 393
rect -381 299 -345 355
rect -289 299 -134 355
rect -78 299 78 355
rect 134 299 289 355
rect 345 299 381 355
rect -381 137 381 299
rect -381 81 -345 137
rect -289 81 -134 137
rect -78 81 78 137
rect 134 81 289 137
rect 345 81 381 137
rect -381 -81 381 81
rect -381 -137 -345 -81
rect -289 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 289 -81
rect 345 -137 381 -81
rect -381 -299 381 -137
rect -381 -355 -345 -299
rect -289 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 289 -299
rect 345 -355 381 -299
rect -381 -393 381 -355
<< via2 >>
rect -345 299 -289 355
rect -134 299 -78 355
rect 78 299 134 355
rect 289 299 345 355
rect -345 81 -289 137
rect -134 81 -78 137
rect 78 81 134 137
rect 289 81 345 137
rect -345 -137 -289 -81
rect -134 -137 -78 -81
rect 78 -137 134 -81
rect 289 -137 345 -81
rect -345 -355 -289 -299
rect -134 -355 -78 -299
rect 78 -355 134 -299
rect 289 -355 345 -299
<< metal3 >>
rect -381 355 381 393
rect -381 299 -345 355
rect -289 299 -134 355
rect -78 299 78 355
rect 134 299 289 355
rect 345 299 381 355
rect -381 137 381 299
rect -381 81 -345 137
rect -289 81 -134 137
rect -78 81 78 137
rect 134 81 289 137
rect 345 81 381 137
rect -381 -81 381 81
rect -381 -137 -345 -81
rect -289 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 289 -81
rect 345 -137 381 -81
rect -381 -299 381 -137
rect -381 -355 -345 -299
rect -289 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 289 -299
rect 345 -355 381 -299
rect -381 -393 381 -355
<< properties >>
string GDS_END 1519734
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1518578
<< end >>
