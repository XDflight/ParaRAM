magic
tech gf180mcuB
timestamp 1666464484
<< properties >>
string GDS_END 1791060
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1790352
<< end >>
