magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 4041
<< polysilicon >>
rect -31 3900 88 3973
rect -31 -74 88 0
use pmos_5p04310590548795_128x8m81  pmos_5p04310590548795_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 4020
<< properties >>
string GDS_END 1120084
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1119770
<< end >>
