magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 568 -141
<< polysilicon >>
rect -31 228 89 300
rect 193 228 313 300
rect -31 -74 89 0
rect 193 -74 313 0
use pmos_5p0431059130203_512x8m81  pmos_5p0431059130203_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 552 348
<< properties >>
string GDS_END 260760
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 260318
<< end >>
