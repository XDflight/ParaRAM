magic
tech gf180mcuB
magscale 1 10
timestamp 1667403392
<< checkpaint >>
rect -2000 -2000 2001 2001
<< end >>
