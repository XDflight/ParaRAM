magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 1120 844
rect 69 506 115 724
rect 244 439 312 676
rect 117 337 312 439
rect 358 337 426 676
rect 582 337 650 676
rect 806 337 874 676
rect 922 476 981 676
rect 922 261 982 476
rect 251 214 982 261
rect 49 60 95 168
rect 251 106 330 214
rect 497 60 543 168
rect 701 106 778 214
rect 945 60 991 168
rect 0 -60 1120 60
<< labels >>
rlabel metal1 s 806 337 874 676 6 A1
port 1 nsew default input
rlabel metal1 s 582 337 650 676 6 A2
port 2 nsew default input
rlabel metal1 s 358 337 426 676 6 A3
port 3 nsew default input
rlabel metal1 s 244 439 312 676 6 A4
port 4 nsew default input
rlabel metal1 s 117 337 312 439 6 A4
port 4 nsew default input
rlabel metal1 s 922 476 981 676 6 ZN
port 5 nsew default output
rlabel metal1 s 922 261 982 476 6 ZN
port 5 nsew default output
rlabel metal1 s 251 214 982 261 6 ZN
port 5 nsew default output
rlabel metal1 s 701 106 778 214 6 ZN
port 5 nsew default output
rlabel metal1 s 251 106 330 214 6 ZN
port 5 nsew default output
rlabel metal1 s 0 724 1120 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 506 115 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 945 60 991 168 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 168 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 168 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1120 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 749006
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 745840
<< end >>
