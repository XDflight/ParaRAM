magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 0 19070 613 24332
rect 286 12610 676 15164
rect 509 10562 1267 11016
rect 488 9531 1373 10562
rect 519 9530 1373 9531
rect 523 3317 1377 5868
rect 392 2240 1377 2696
<< psubdiff >>
rect 707 8816 1183 8876
rect 707 8770 764 8816
rect 810 8770 922 8816
rect 968 8770 1080 8816
rect 1126 8770 1183 8816
rect 707 8710 1183 8770
<< nsubdiff >>
rect 652 10811 1124 10868
rect 652 10765 707 10811
rect 753 10765 865 10811
rect 911 10765 1023 10811
rect 1069 10765 1124 10811
rect 652 10708 1124 10765
rect 535 2491 690 2548
rect 535 2445 589 2491
rect 635 2445 690 2491
rect 535 2388 690 2445
rect 1079 2491 1234 2548
rect 1079 2445 1133 2491
rect 1179 2445 1234 2491
rect 1079 2388 1234 2445
<< psubdiffcont >>
rect 764 8770 810 8816
rect 922 8770 968 8816
rect 1080 8770 1126 8816
<< nsubdiffcont >>
rect 707 10765 753 10811
rect 865 10765 911 10811
rect 1023 10765 1069 10811
rect 589 2445 635 2491
rect 1133 2445 1179 2491
<< polysilicon >>
rect 795 9629 872 9671
rect 1019 9629 1096 9671
rect 774 9612 894 9629
rect 998 9612 1118 9629
rect 774 9596 1118 9612
rect 774 9550 1407 9596
rect 774 9504 1129 9550
rect 1175 9504 1287 9550
rect 1333 9504 1407 9550
rect 774 9458 1407 9504
rect 774 9449 1118 9458
rect 774 9388 894 9449
rect 998 9388 1118 9449
rect 774 9009 894 9091
rect 998 9009 1118 9091
rect 778 5944 898 6006
rect 1002 5944 1122 6006
rect 778 5935 1122 5944
rect 471 5889 1122 5935
rect 471 5843 545 5889
rect 591 5843 703 5889
rect 749 5843 1122 5889
rect 471 5797 1122 5843
rect 778 5786 1122 5797
rect 778 5770 898 5786
rect 1002 5770 1122 5786
rect 799 5727 876 5770
rect 1023 5727 1100 5770
<< polycontact >>
rect 1129 9504 1175 9550
rect 1287 9504 1333 9550
rect 545 5843 591 5889
rect 703 5843 749 5889
<< metal1 >>
rect 808 19210 1022 20572
rect 310 13516 869 13636
rect 310 11789 426 13516
rect 1049 13117 1291 13414
rect 310 11669 1441 11789
rect 672 10811 1104 10848
rect 672 10765 707 10811
rect 753 10765 865 10811
rect 911 10765 1023 10811
rect 1069 10765 1104 10811
rect 672 10728 1104 10765
rect 887 9601 1004 9986
rect 486 9526 1004 9601
rect 1324 9587 1441 11669
rect 486 5926 558 9526
rect 887 9263 1004 9526
rect 1094 9550 1441 9587
rect 1094 9504 1129 9550
rect 1175 9504 1287 9550
rect 1333 9504 1441 9550
rect 1094 9467 1441 9504
rect 663 8867 780 9141
rect 1111 8867 1228 9141
rect 663 8816 1228 8867
rect 663 8770 764 8816
rect 810 8770 922 8816
rect 968 8770 1080 8816
rect 1126 8770 1228 8816
rect 663 8719 1228 8770
rect 663 6922 780 8719
rect 486 5889 784 5926
rect 486 5843 545 5889
rect 591 5843 703 5889
rect 749 5843 784 5889
rect 486 5806 784 5843
rect 892 5580 1008 6967
rect 1111 6922 1228 8719
rect 668 2528 784 3722
rect 1116 2528 1232 3722
rect 555 2491 784 2528
rect 555 2445 589 2491
rect 635 2445 784 2491
rect 555 2408 784 2445
rect 887 2245 1017 2512
rect 1099 2491 1232 2528
rect 1099 2445 1133 2491
rect 1179 2445 1232 2491
rect 1099 2408 1232 2445
rect 839 0 1061 2245
<< metal2 >>
rect 728 24553 848 24714
rect 685 24455 848 24553
rect 1028 24553 1148 24714
rect 1028 24455 1156 24553
rect 685 24160 741 24455
rect 1100 24160 1156 24455
rect 887 0 1017 7812
<< metal3 >>
rect 167 22500 1737 24309
rect 222 16619 1737 18618
rect 117 16293 1737 16508
rect 117 15971 1737 16187
rect 117 15650 1737 15865
rect 117 15328 1737 15543
rect 117 14636 1447 14851
rect 117 14314 1447 14529
rect 117 13992 1447 14207
rect 117 13670 1447 13886
rect 222 13122 1737 13564
rect 222 12011 1737 12466
rect 264 8200 1241 10923
rect 264 4512 1241 7914
rect 189 3646 1241 4363
rect 189 2220 1241 3031
rect 264 359 889 1675
use M1_NWELL$$44998700_256x8m81_0  M1_NWELL$$44998700_256x8m81_0_0
timestamp 1666464484
transform 1 0 1156 0 1 2468
box 0 0 1 1
use M1_NWELL$$44998700_256x8m81_0  M1_NWELL$$44998700_256x8m81_0_1
timestamp 1666464484
transform 1 0 612 0 1 2468
box 0 0 1 1
use M1_NWELL$$46277676_256x8m81_0  M1_NWELL$$46277676_256x8m81_0_0
timestamp 1666464484
transform 1 0 888 0 1 10788
box 0 0 1 1
use M1_POLY2$$46559276_256x8m81  M1_POLY2$$46559276_256x8m81_0
timestamp 1666464484
transform -1 0 647 0 1 5866
box 0 0 1 1
use M1_POLY2$$46559276_256x8m81  M1_POLY2$$46559276_256x8m81_1
timestamp 1666464484
transform 1 0 1231 0 1 9527
box 0 0 1 1
use M1_PSUB$$46274604_256x8m81  M1_PSUB$$46274604_256x8m81_0
timestamp 1666464484
transform 1 0 945 0 1 8793
box 0 0 1 1
use M2_M1$$47117356_256x8m81  M2_M1$$47117356_256x8m81_0
timestamp 1666464484
transform 1 0 952 0 1 5141
box -65 -2678 65 2678
use nmos_5p04310590878154_256x8m81  nmos_5p04310590878154_256x8m81_0
timestamp 1666464484
transform 1 0 778 0 1 6007
box -88 -44 432 1744
use nmos_5p04310590878156_256x8m81  nmos_5p04310590878156_256x8m81_0
timestamp 1666464484
transform 1 0 774 0 1 9092
box -88 -44 432 320
use pmos_5p04310590878153_256x8m81  pmos_5p04310590878153_256x8m81_0
timestamp 1666464484
transform 1 0 774 0 1 9672
box -208 -120 552 822
use pmos_5p04310590878155_256x8m81  pmos_5p04310590878155_256x8m81_0
timestamp 1666464484
transform 1 0 778 0 -1 5726
box -208 -120 552 2248
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_0
timestamp 1666464484
transform 1 0 680 0 1 7501
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_1
timestamp 1666464484
transform 1 0 680 0 1 6358
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_2
timestamp 1666464484
transform 1 0 680 0 1 6963
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_3
timestamp 1666464484
transform 1 0 684 0 1 2513
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_4
timestamp 1666464484
transform 1 0 684 0 1 2699
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_5
timestamp 1666464484
transform 1 0 1121 0 1 7501
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_6
timestamp 1666464484
transform 1 0 1121 0 1 6358
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_7
timestamp 1666464484
transform 1 0 1121 0 1 6963
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_8
timestamp 1666464484
transform 1 0 1123 0 1 9940
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_9
timestamp 1666464484
transform 1 0 1126 0 1 2699
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_10
timestamp 1666464484
transform 1 0 1126 0 1 2513
box 0 -1 93 308
use via1_2_x2_256x8m81_0  via1_2_x2_256x8m81_0_11
timestamp 1666464484
transform 1 0 675 0 1 9940
box 0 -1 93 308
use via1_2_x2_R90_256x8m81_0  via1_2_x2_R90_256x8m81_0_0
timestamp 1666464484
transform 0 -1 1025 1 0 10740
box 0 -1 93 308
use via1_2_x2_R270_256x8m81_0  via1_2_x2_R270_256x8m81_0_0
timestamp 1666464484
transform 0 1 632 -1 0 13408
box -1 -1 96 308
use ypass_gate_256x8m81_0  ypass_gate_256x8m81_0_0
timestamp 1666464484
transform -1 0 1233 0 1 11962
box -221 -1 930 12370
<< labels >>
rlabel metal1 s 877 8804 877 8804 4 vss
port 1 nsew
rlabel metal1 s 875 22284 875 22284 4 pcb
port 2 nsew
rlabel metal1 s 875 22284 875 22284 4 pcb
port 2 nsew
rlabel metal1 s 965 158 965 158 4 tblhl
port 3 nsew
rlabel metal3 s 379 18693 379 18693 4 vss
port 1 nsew
rlabel metal3 s 379 24134 379 24134 4 vdd
port 4 nsew
rlabel metal3 s 379 13372 379 13372 4 vdd
port 4 nsew
rlabel metal3 s 379 10706 379 10706 4 vdd
port 4 nsew
rlabel metal3 s 379 4225 379 4225 4 vdd
port 4 nsew
rlabel metal3 s 482 12248 482 12248 4 vss
port 1 nsew
<< properties >>
string GDS_END 853284
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 847500
<< end >>
