magic
tech gf180mcuA
magscale 1 10
timestamp 1667403433
<< checkpaint >>
rect -2000 -2000 2001 2001
<< end >>
