magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -2449 102 2449 159
rect -2449 56 -2390 102
rect -2344 56 -2227 102
rect -2181 56 -2064 102
rect -2018 56 -1900 102
rect -1854 56 -1737 102
rect -1691 56 -1574 102
rect -1528 56 -1411 102
rect -1365 56 -1247 102
rect -1201 56 -1084 102
rect -1038 56 -921 102
rect -875 56 -758 102
rect -712 56 -595 102
rect -549 56 -431 102
rect -385 56 -268 102
rect -222 56 -105 102
rect -59 56 59 102
rect 105 56 222 102
rect 268 56 385 102
rect 431 56 549 102
rect 595 56 712 102
rect 758 56 875 102
rect 921 56 1038 102
rect 1084 56 1201 102
rect 1247 56 1365 102
rect 1411 56 1528 102
rect 1574 56 1691 102
rect 1737 56 1854 102
rect 1900 56 2018 102
rect 2064 56 2181 102
rect 2227 56 2344 102
rect 2390 56 2449 102
rect -2449 -56 2449 56
rect -2449 -102 -2390 -56
rect -2344 -102 -2227 -56
rect -2181 -102 -2064 -56
rect -2018 -102 -1900 -56
rect -1854 -102 -1737 -56
rect -1691 -102 -1574 -56
rect -1528 -102 -1411 -56
rect -1365 -102 -1247 -56
rect -1201 -102 -1084 -56
rect -1038 -102 -921 -56
rect -875 -102 -758 -56
rect -712 -102 -595 -56
rect -549 -102 -431 -56
rect -385 -102 -268 -56
rect -222 -102 -105 -56
rect -59 -102 59 -56
rect 105 -102 222 -56
rect 268 -102 385 -56
rect 431 -102 549 -56
rect 595 -102 712 -56
rect 758 -102 875 -56
rect 921 -102 1038 -56
rect 1084 -102 1201 -56
rect 1247 -102 1365 -56
rect 1411 -102 1528 -56
rect 1574 -102 1691 -56
rect 1737 -102 1854 -56
rect 1900 -102 2018 -56
rect 2064 -102 2181 -56
rect 2227 -102 2344 -56
rect 2390 -102 2449 -56
rect -2449 -159 2449 -102
<< psubdiffcont >>
rect -2390 56 -2344 102
rect -2227 56 -2181 102
rect -2064 56 -2018 102
rect -1900 56 -1854 102
rect -1737 56 -1691 102
rect -1574 56 -1528 102
rect -1411 56 -1365 102
rect -1247 56 -1201 102
rect -1084 56 -1038 102
rect -921 56 -875 102
rect -758 56 -712 102
rect -595 56 -549 102
rect -431 56 -385 102
rect -268 56 -222 102
rect -105 56 -59 102
rect 59 56 105 102
rect 222 56 268 102
rect 385 56 431 102
rect 549 56 595 102
rect 712 56 758 102
rect 875 56 921 102
rect 1038 56 1084 102
rect 1201 56 1247 102
rect 1365 56 1411 102
rect 1528 56 1574 102
rect 1691 56 1737 102
rect 1854 56 1900 102
rect 2018 56 2064 102
rect 2181 56 2227 102
rect 2344 56 2390 102
rect -2390 -102 -2344 -56
rect -2227 -102 -2181 -56
rect -2064 -102 -2018 -56
rect -1900 -102 -1854 -56
rect -1737 -102 -1691 -56
rect -1574 -102 -1528 -56
rect -1411 -102 -1365 -56
rect -1247 -102 -1201 -56
rect -1084 -102 -1038 -56
rect -921 -102 -875 -56
rect -758 -102 -712 -56
rect -595 -102 -549 -56
rect -431 -102 -385 -56
rect -268 -102 -222 -56
rect -105 -102 -59 -56
rect 59 -102 105 -56
rect 222 -102 268 -56
rect 385 -102 431 -56
rect 549 -102 595 -56
rect 712 -102 758 -56
rect 875 -102 921 -56
rect 1038 -102 1084 -56
rect 1201 -102 1247 -56
rect 1365 -102 1411 -56
rect 1528 -102 1574 -56
rect 1691 -102 1737 -56
rect 1854 -102 1900 -56
rect 2018 -102 2064 -56
rect 2181 -102 2227 -56
rect 2344 -102 2390 -56
<< metal1 >>
rect -2440 102 2440 150
rect -2440 56 -2390 102
rect -2344 56 -2227 102
rect -2181 56 -2064 102
rect -2018 56 -1900 102
rect -1854 56 -1737 102
rect -1691 56 -1574 102
rect -1528 56 -1411 102
rect -1365 56 -1247 102
rect -1201 56 -1084 102
rect -1038 56 -921 102
rect -875 56 -758 102
rect -712 56 -595 102
rect -549 56 -431 102
rect -385 56 -268 102
rect -222 56 -105 102
rect -59 56 59 102
rect 105 56 222 102
rect 268 56 385 102
rect 431 56 549 102
rect 595 56 712 102
rect 758 56 875 102
rect 921 56 1038 102
rect 1084 56 1201 102
rect 1247 56 1365 102
rect 1411 56 1528 102
rect 1574 56 1691 102
rect 1737 56 1854 102
rect 1900 56 2018 102
rect 2064 56 2181 102
rect 2227 56 2344 102
rect 2390 56 2440 102
rect -2440 -56 2440 56
rect -2440 -102 -2390 -56
rect -2344 -102 -2227 -56
rect -2181 -102 -2064 -56
rect -2018 -102 -1900 -56
rect -1854 -102 -1737 -56
rect -1691 -102 -1574 -56
rect -1528 -102 -1411 -56
rect -1365 -102 -1247 -56
rect -1201 -102 -1084 -56
rect -1038 -102 -921 -56
rect -875 -102 -758 -56
rect -712 -102 -595 -56
rect -549 -102 -431 -56
rect -385 -102 -268 -56
rect -222 -102 -105 -56
rect -59 -102 59 -56
rect 105 -102 222 -56
rect 268 -102 385 -56
rect 431 -102 549 -56
rect 595 -102 712 -56
rect 758 -102 875 -56
rect 921 -102 1038 -56
rect 1084 -102 1201 -56
rect 1247 -102 1365 -56
rect 1411 -102 1528 -56
rect 1574 -102 1691 -56
rect 1737 -102 1854 -56
rect 1900 -102 2018 -56
rect 2064 -102 2181 -56
rect 2227 -102 2344 -56
rect 2390 -102 2440 -56
rect -2440 -150 2440 -102
<< properties >>
string GDS_END 830028
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 825992
<< end >>
