magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -143 75 143 81
rect -143 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 143 75
rect -143 13 143 49
rect -143 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 143 13
rect -143 -49 143 -13
rect -143 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 143 -49
rect -143 -81 143 -75
<< via1 >>
rect -137 49 -111 75
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect 111 49 137 75
rect -137 -13 -111 13
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect 111 -13 137 13
rect -137 -75 -111 -49
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect 111 -75 137 -49
<< metal2 >>
rect -143 75 143 81
rect -143 49 -137 75
rect -111 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 111 75
rect 137 49 143 75
rect -143 13 143 49
rect -143 -13 -137 13
rect -111 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 111 13
rect 137 -13 143 13
rect -143 -49 143 -13
rect -143 -75 -137 -49
rect -111 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 111 -49
rect 137 -75 143 -49
rect -143 -81 143 -75
<< properties >>
string GDS_END 1908884
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1907792
<< end >>
