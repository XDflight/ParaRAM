magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 395 85602 414
rect -42 349 -23 395
rect 23 349 101 395
rect 147 349 225 395
rect 271 349 349 395
rect 395 349 473 395
rect 519 349 597 395
rect 643 349 721 395
rect 767 349 845 395
rect 891 349 969 395
rect 1015 349 1093 395
rect 1139 349 1217 395
rect 1263 349 1341 395
rect 1387 349 1465 395
rect 1511 349 1589 395
rect 1635 349 1713 395
rect 1759 349 1837 395
rect 1883 349 1961 395
rect 2007 349 2085 395
rect 2131 349 2209 395
rect 2255 349 2333 395
rect 2379 349 2457 395
rect 2503 349 2581 395
rect 2627 349 2705 395
rect 2751 349 2829 395
rect 2875 349 2953 395
rect 2999 349 3077 395
rect 3123 349 3201 395
rect 3247 349 3325 395
rect 3371 349 3449 395
rect 3495 349 3573 395
rect 3619 349 3697 395
rect 3743 349 3821 395
rect 3867 349 3945 395
rect 3991 349 4069 395
rect 4115 349 4193 395
rect 4239 349 4317 395
rect 4363 349 4441 395
rect 4487 349 4565 395
rect 4611 349 4689 395
rect 4735 349 4813 395
rect 4859 349 4937 395
rect 4983 349 5061 395
rect 5107 349 5185 395
rect 5231 349 5309 395
rect 5355 349 5433 395
rect 5479 349 5557 395
rect 5603 349 5681 395
rect 5727 349 5805 395
rect 5851 349 5929 395
rect 5975 349 6053 395
rect 6099 349 6177 395
rect 6223 349 6301 395
rect 6347 349 6425 395
rect 6471 349 6549 395
rect 6595 349 6673 395
rect 6719 349 6797 395
rect 6843 349 6921 395
rect 6967 349 7045 395
rect 7091 349 7169 395
rect 7215 349 7293 395
rect 7339 349 7417 395
rect 7463 349 7541 395
rect 7587 349 7665 395
rect 7711 349 7789 395
rect 7835 349 7913 395
rect 7959 349 8037 395
rect 8083 349 8161 395
rect 8207 349 8285 395
rect 8331 349 8409 395
rect 8455 349 8533 395
rect 8579 349 8657 395
rect 8703 349 8781 395
rect 8827 349 8905 395
rect 8951 349 9029 395
rect 9075 349 9153 395
rect 9199 349 9277 395
rect 9323 349 9401 395
rect 9447 349 9525 395
rect 9571 349 9649 395
rect 9695 349 9773 395
rect 9819 349 9897 395
rect 9943 349 10021 395
rect 10067 349 10145 395
rect 10191 349 10269 395
rect 10315 349 10393 395
rect 10439 349 10517 395
rect 10563 349 10641 395
rect 10687 349 10765 395
rect 10811 349 10889 395
rect 10935 349 11013 395
rect 11059 349 11137 395
rect 11183 349 11261 395
rect 11307 349 11385 395
rect 11431 349 11509 395
rect 11555 349 11633 395
rect 11679 349 11757 395
rect 11803 349 11881 395
rect 11927 349 12005 395
rect 12051 349 12129 395
rect 12175 349 12253 395
rect 12299 349 12377 395
rect 12423 349 12501 395
rect 12547 349 12625 395
rect 12671 349 12749 395
rect 12795 349 12873 395
rect 12919 349 12997 395
rect 13043 349 13121 395
rect 13167 349 13245 395
rect 13291 349 13369 395
rect 13415 349 13493 395
rect 13539 349 13617 395
rect 13663 349 13741 395
rect 13787 349 13865 395
rect 13911 349 13989 395
rect 14035 349 14113 395
rect 14159 349 14237 395
rect 14283 349 14361 395
rect 14407 349 14485 395
rect 14531 349 14609 395
rect 14655 349 14733 395
rect 14779 349 14857 395
rect 14903 349 14981 395
rect 15027 349 15105 395
rect 15151 349 15229 395
rect 15275 349 15353 395
rect 15399 349 15477 395
rect 15523 349 15601 395
rect 15647 349 15725 395
rect 15771 349 15849 395
rect 15895 349 15973 395
rect 16019 349 16097 395
rect 16143 349 16221 395
rect 16267 349 16345 395
rect 16391 349 16469 395
rect 16515 349 16593 395
rect 16639 349 16717 395
rect 16763 349 16841 395
rect 16887 349 16965 395
rect 17011 349 17089 395
rect 17135 349 17213 395
rect 17259 349 17337 395
rect 17383 349 17461 395
rect 17507 349 17585 395
rect 17631 349 17709 395
rect 17755 349 17833 395
rect 17879 349 17957 395
rect 18003 349 18081 395
rect 18127 349 18205 395
rect 18251 349 18329 395
rect 18375 349 18453 395
rect 18499 349 18577 395
rect 18623 349 18701 395
rect 18747 349 18825 395
rect 18871 349 18949 395
rect 18995 349 19073 395
rect 19119 349 19197 395
rect 19243 349 19321 395
rect 19367 349 19445 395
rect 19491 349 19569 395
rect 19615 349 19693 395
rect 19739 349 19817 395
rect 19863 349 19941 395
rect 19987 349 20065 395
rect 20111 349 20189 395
rect 20235 349 20313 395
rect 20359 349 20437 395
rect 20483 349 20561 395
rect 20607 349 20685 395
rect 20731 349 20809 395
rect 20855 349 20933 395
rect 20979 349 21057 395
rect 21103 349 21181 395
rect 21227 349 21305 395
rect 21351 349 21429 395
rect 21475 349 21553 395
rect 21599 349 21677 395
rect 21723 349 21801 395
rect 21847 349 21925 395
rect 21971 349 22049 395
rect 22095 349 22173 395
rect 22219 349 22297 395
rect 22343 349 22421 395
rect 22467 349 22545 395
rect 22591 349 22669 395
rect 22715 349 22793 395
rect 22839 349 22917 395
rect 22963 349 23041 395
rect 23087 349 23165 395
rect 23211 349 23289 395
rect 23335 349 23413 395
rect 23459 349 23537 395
rect 23583 349 23661 395
rect 23707 349 23785 395
rect 23831 349 23909 395
rect 23955 349 24033 395
rect 24079 349 24157 395
rect 24203 349 24281 395
rect 24327 349 24405 395
rect 24451 349 24529 395
rect 24575 349 24653 395
rect 24699 349 24777 395
rect 24823 349 24901 395
rect 24947 349 25025 395
rect 25071 349 25149 395
rect 25195 349 25273 395
rect 25319 349 25397 395
rect 25443 349 25521 395
rect 25567 349 25645 395
rect 25691 349 25769 395
rect 25815 349 25893 395
rect 25939 349 26017 395
rect 26063 349 26141 395
rect 26187 349 26265 395
rect 26311 349 26389 395
rect 26435 349 26513 395
rect 26559 349 26637 395
rect 26683 349 26761 395
rect 26807 349 26885 395
rect 26931 349 27009 395
rect 27055 349 27133 395
rect 27179 349 27257 395
rect 27303 349 27381 395
rect 27427 349 27505 395
rect 27551 349 27629 395
rect 27675 349 27753 395
rect 27799 349 27877 395
rect 27923 349 28001 395
rect 28047 349 28125 395
rect 28171 349 28249 395
rect 28295 349 28373 395
rect 28419 349 28497 395
rect 28543 349 28621 395
rect 28667 349 28745 395
rect 28791 349 28869 395
rect 28915 349 28993 395
rect 29039 349 29117 395
rect 29163 349 29241 395
rect 29287 349 29365 395
rect 29411 349 29489 395
rect 29535 349 29613 395
rect 29659 349 29737 395
rect 29783 349 29861 395
rect 29907 349 29985 395
rect 30031 349 30109 395
rect 30155 349 30233 395
rect 30279 349 30357 395
rect 30403 349 30481 395
rect 30527 349 30605 395
rect 30651 349 30729 395
rect 30775 349 30853 395
rect 30899 349 30977 395
rect 31023 349 31101 395
rect 31147 349 31225 395
rect 31271 349 31349 395
rect 31395 349 31473 395
rect 31519 349 31597 395
rect 31643 349 31721 395
rect 31767 349 31845 395
rect 31891 349 31969 395
rect 32015 349 32093 395
rect 32139 349 32217 395
rect 32263 349 32341 395
rect 32387 349 32465 395
rect 32511 349 32589 395
rect 32635 349 32713 395
rect 32759 349 32837 395
rect 32883 349 32961 395
rect 33007 349 33085 395
rect 33131 349 33209 395
rect 33255 349 33333 395
rect 33379 349 33457 395
rect 33503 349 33581 395
rect 33627 349 33705 395
rect 33751 349 33829 395
rect 33875 349 33953 395
rect 33999 349 34077 395
rect 34123 349 34201 395
rect 34247 349 34325 395
rect 34371 349 34449 395
rect 34495 349 34573 395
rect 34619 349 34697 395
rect 34743 349 34821 395
rect 34867 349 34945 395
rect 34991 349 35069 395
rect 35115 349 35193 395
rect 35239 349 35317 395
rect 35363 349 35441 395
rect 35487 349 35565 395
rect 35611 349 35689 395
rect 35735 349 35813 395
rect 35859 349 35937 395
rect 35983 349 36061 395
rect 36107 349 36185 395
rect 36231 349 36309 395
rect 36355 349 36433 395
rect 36479 349 36557 395
rect 36603 349 36681 395
rect 36727 349 36805 395
rect 36851 349 36929 395
rect 36975 349 37053 395
rect 37099 349 37177 395
rect 37223 349 37301 395
rect 37347 349 37425 395
rect 37471 349 37549 395
rect 37595 349 37673 395
rect 37719 349 37797 395
rect 37843 349 37921 395
rect 37967 349 38045 395
rect 38091 349 38169 395
rect 38215 349 38293 395
rect 38339 349 38417 395
rect 38463 349 38541 395
rect 38587 349 38665 395
rect 38711 349 38789 395
rect 38835 349 38913 395
rect 38959 349 39037 395
rect 39083 349 39161 395
rect 39207 349 39285 395
rect 39331 349 39409 395
rect 39455 349 39533 395
rect 39579 349 39657 395
rect 39703 349 39781 395
rect 39827 349 39905 395
rect 39951 349 40029 395
rect 40075 349 40153 395
rect 40199 349 40277 395
rect 40323 349 40401 395
rect 40447 349 40525 395
rect 40571 349 40649 395
rect 40695 349 40773 395
rect 40819 349 40897 395
rect 40943 349 41021 395
rect 41067 349 41145 395
rect 41191 349 41269 395
rect 41315 349 41393 395
rect 41439 349 41517 395
rect 41563 349 41641 395
rect 41687 349 41765 395
rect 41811 349 41889 395
rect 41935 349 42013 395
rect 42059 349 42137 395
rect 42183 349 42261 395
rect 42307 349 42385 395
rect 42431 349 42509 395
rect 42555 349 42633 395
rect 42679 349 42757 395
rect 42803 349 42881 395
rect 42927 349 43005 395
rect 43051 349 43129 395
rect 43175 349 43253 395
rect 43299 349 43377 395
rect 43423 349 43501 395
rect 43547 349 43625 395
rect 43671 349 43749 395
rect 43795 349 43873 395
rect 43919 349 43997 395
rect 44043 349 44121 395
rect 44167 349 44245 395
rect 44291 349 44369 395
rect 44415 349 44493 395
rect 44539 349 44617 395
rect 44663 349 44741 395
rect 44787 349 44865 395
rect 44911 349 44989 395
rect 45035 349 45113 395
rect 45159 349 45237 395
rect 45283 349 45361 395
rect 45407 349 45485 395
rect 45531 349 45609 395
rect 45655 349 45733 395
rect 45779 349 45857 395
rect 45903 349 45981 395
rect 46027 349 46105 395
rect 46151 349 46229 395
rect 46275 349 46353 395
rect 46399 349 46477 395
rect 46523 349 46601 395
rect 46647 349 46725 395
rect 46771 349 46849 395
rect 46895 349 46973 395
rect 47019 349 47097 395
rect 47143 349 47221 395
rect 47267 349 47345 395
rect 47391 349 47469 395
rect 47515 349 47593 395
rect 47639 349 47717 395
rect 47763 349 47841 395
rect 47887 349 47965 395
rect 48011 349 48089 395
rect 48135 349 48213 395
rect 48259 349 48337 395
rect 48383 349 48461 395
rect 48507 349 48585 395
rect 48631 349 48709 395
rect 48755 349 48833 395
rect 48879 349 48957 395
rect 49003 349 49081 395
rect 49127 349 49205 395
rect 49251 349 49329 395
rect 49375 349 49453 395
rect 49499 349 49577 395
rect 49623 349 49701 395
rect 49747 349 49825 395
rect 49871 349 49949 395
rect 49995 349 50073 395
rect 50119 349 50197 395
rect 50243 349 50321 395
rect 50367 349 50445 395
rect 50491 349 50569 395
rect 50615 349 50693 395
rect 50739 349 50817 395
rect 50863 349 50941 395
rect 50987 349 51065 395
rect 51111 349 51189 395
rect 51235 349 51313 395
rect 51359 349 51437 395
rect 51483 349 51561 395
rect 51607 349 51685 395
rect 51731 349 51809 395
rect 51855 349 51933 395
rect 51979 349 52057 395
rect 52103 349 52181 395
rect 52227 349 52305 395
rect 52351 349 52429 395
rect 52475 349 52553 395
rect 52599 349 52677 395
rect 52723 349 52801 395
rect 52847 349 52925 395
rect 52971 349 53049 395
rect 53095 349 53173 395
rect 53219 349 53297 395
rect 53343 349 53421 395
rect 53467 349 53545 395
rect 53591 349 53669 395
rect 53715 349 53793 395
rect 53839 349 53917 395
rect 53963 349 54041 395
rect 54087 349 54165 395
rect 54211 349 54289 395
rect 54335 349 54413 395
rect 54459 349 54537 395
rect 54583 349 54661 395
rect 54707 349 54785 395
rect 54831 349 54909 395
rect 54955 349 55033 395
rect 55079 349 55157 395
rect 55203 349 55281 395
rect 55327 349 55405 395
rect 55451 349 55529 395
rect 55575 349 55653 395
rect 55699 349 55777 395
rect 55823 349 55901 395
rect 55947 349 56025 395
rect 56071 349 56149 395
rect 56195 349 56273 395
rect 56319 349 56397 395
rect 56443 349 56521 395
rect 56567 349 56645 395
rect 56691 349 56769 395
rect 56815 349 56893 395
rect 56939 349 57017 395
rect 57063 349 57141 395
rect 57187 349 57265 395
rect 57311 349 57389 395
rect 57435 349 57513 395
rect 57559 349 57637 395
rect 57683 349 57761 395
rect 57807 349 57885 395
rect 57931 349 58009 395
rect 58055 349 58133 395
rect 58179 349 58257 395
rect 58303 349 58381 395
rect 58427 349 58505 395
rect 58551 349 58629 395
rect 58675 349 58753 395
rect 58799 349 58877 395
rect 58923 349 59001 395
rect 59047 349 59125 395
rect 59171 349 59249 395
rect 59295 349 59373 395
rect 59419 349 59497 395
rect 59543 349 59621 395
rect 59667 349 59745 395
rect 59791 349 59869 395
rect 59915 349 59993 395
rect 60039 349 60117 395
rect 60163 349 60241 395
rect 60287 349 60365 395
rect 60411 349 60489 395
rect 60535 349 60613 395
rect 60659 349 60737 395
rect 60783 349 60861 395
rect 60907 349 60985 395
rect 61031 349 61109 395
rect 61155 349 61233 395
rect 61279 349 61357 395
rect 61403 349 61481 395
rect 61527 349 61605 395
rect 61651 349 61729 395
rect 61775 349 61853 395
rect 61899 349 61977 395
rect 62023 349 62101 395
rect 62147 349 62225 395
rect 62271 349 62349 395
rect 62395 349 62473 395
rect 62519 349 62597 395
rect 62643 349 62721 395
rect 62767 349 62845 395
rect 62891 349 62969 395
rect 63015 349 63093 395
rect 63139 349 63217 395
rect 63263 349 63341 395
rect 63387 349 63465 395
rect 63511 349 63589 395
rect 63635 349 63713 395
rect 63759 349 63837 395
rect 63883 349 63961 395
rect 64007 349 64085 395
rect 64131 349 64209 395
rect 64255 349 64333 395
rect 64379 349 64457 395
rect 64503 349 64581 395
rect 64627 349 64705 395
rect 64751 349 64829 395
rect 64875 349 64953 395
rect 64999 349 65077 395
rect 65123 349 65201 395
rect 65247 349 65325 395
rect 65371 349 65449 395
rect 65495 349 65573 395
rect 65619 349 65697 395
rect 65743 349 65821 395
rect 65867 349 65945 395
rect 65991 349 66069 395
rect 66115 349 66193 395
rect 66239 349 66317 395
rect 66363 349 66441 395
rect 66487 349 66565 395
rect 66611 349 66689 395
rect 66735 349 66813 395
rect 66859 349 66937 395
rect 66983 349 67061 395
rect 67107 349 67185 395
rect 67231 349 67309 395
rect 67355 349 67433 395
rect 67479 349 67557 395
rect 67603 349 67681 395
rect 67727 349 67805 395
rect 67851 349 67929 395
rect 67975 349 68053 395
rect 68099 349 68177 395
rect 68223 349 68301 395
rect 68347 349 68425 395
rect 68471 349 68549 395
rect 68595 349 68673 395
rect 68719 349 68797 395
rect 68843 349 68921 395
rect 68967 349 69045 395
rect 69091 349 69169 395
rect 69215 349 69293 395
rect 69339 349 69417 395
rect 69463 349 69541 395
rect 69587 349 69665 395
rect 69711 349 69789 395
rect 69835 349 69913 395
rect 69959 349 70037 395
rect 70083 349 70161 395
rect 70207 349 70285 395
rect 70331 349 70409 395
rect 70455 349 70533 395
rect 70579 349 70657 395
rect 70703 349 70781 395
rect 70827 349 70905 395
rect 70951 349 71029 395
rect 71075 349 71153 395
rect 71199 349 71277 395
rect 71323 349 71401 395
rect 71447 349 71525 395
rect 71571 349 71649 395
rect 71695 349 71773 395
rect 71819 349 71897 395
rect 71943 349 72021 395
rect 72067 349 72145 395
rect 72191 349 72269 395
rect 72315 349 72393 395
rect 72439 349 72517 395
rect 72563 349 72641 395
rect 72687 349 72765 395
rect 72811 349 72889 395
rect 72935 349 73013 395
rect 73059 349 73137 395
rect 73183 349 73261 395
rect 73307 349 73385 395
rect 73431 349 73509 395
rect 73555 349 73633 395
rect 73679 349 73757 395
rect 73803 349 73881 395
rect 73927 349 74005 395
rect 74051 349 74129 395
rect 74175 349 74253 395
rect 74299 349 74377 395
rect 74423 349 74501 395
rect 74547 349 74625 395
rect 74671 349 74749 395
rect 74795 349 74873 395
rect 74919 349 74997 395
rect 75043 349 75121 395
rect 75167 349 75245 395
rect 75291 349 75369 395
rect 75415 349 75493 395
rect 75539 349 75617 395
rect 75663 349 75741 395
rect 75787 349 75865 395
rect 75911 349 75989 395
rect 76035 349 76113 395
rect 76159 349 76237 395
rect 76283 349 76361 395
rect 76407 349 76485 395
rect 76531 349 76609 395
rect 76655 349 76733 395
rect 76779 349 76857 395
rect 76903 349 76981 395
rect 77027 349 77105 395
rect 77151 349 77229 395
rect 77275 349 77353 395
rect 77399 349 77477 395
rect 77523 349 77601 395
rect 77647 349 77725 395
rect 77771 349 77849 395
rect 77895 349 77973 395
rect 78019 349 78097 395
rect 78143 349 78221 395
rect 78267 349 78345 395
rect 78391 349 78469 395
rect 78515 349 78593 395
rect 78639 349 78717 395
rect 78763 349 78841 395
rect 78887 349 78965 395
rect 79011 349 79089 395
rect 79135 349 79213 395
rect 79259 349 79337 395
rect 79383 349 79461 395
rect 79507 349 79585 395
rect 79631 349 79709 395
rect 79755 349 79833 395
rect 79879 349 79957 395
rect 80003 349 80081 395
rect 80127 349 80205 395
rect 80251 349 80329 395
rect 80375 349 80453 395
rect 80499 349 80577 395
rect 80623 349 80701 395
rect 80747 349 80825 395
rect 80871 349 80949 395
rect 80995 349 81073 395
rect 81119 349 81197 395
rect 81243 349 81321 395
rect 81367 349 81445 395
rect 81491 349 81569 395
rect 81615 349 81693 395
rect 81739 349 81817 395
rect 81863 349 81941 395
rect 81987 349 82065 395
rect 82111 349 82189 395
rect 82235 349 82313 395
rect 82359 349 82437 395
rect 82483 349 82561 395
rect 82607 349 82685 395
rect 82731 349 82809 395
rect 82855 349 82933 395
rect 82979 349 83057 395
rect 83103 349 83181 395
rect 83227 349 83305 395
rect 83351 349 83429 395
rect 83475 349 83553 395
rect 83599 349 83677 395
rect 83723 349 83801 395
rect 83847 349 83925 395
rect 83971 349 84049 395
rect 84095 349 84173 395
rect 84219 349 84297 395
rect 84343 349 84421 395
rect 84467 349 84545 395
rect 84591 349 84669 395
rect 84715 349 84793 395
rect 84839 349 84917 395
rect 84963 349 85041 395
rect 85087 349 85165 395
rect 85211 349 85289 395
rect 85335 349 85413 395
rect 85459 349 85537 395
rect 85583 349 85602 395
rect -42 271 85602 349
rect -42 225 -23 271
rect 23 225 101 271
rect 147 225 225 271
rect 271 225 349 271
rect 395 225 473 271
rect 519 225 597 271
rect 643 225 721 271
rect 767 225 845 271
rect 891 225 969 271
rect 1015 225 1093 271
rect 1139 225 1217 271
rect 1263 225 1341 271
rect 1387 225 1465 271
rect 1511 225 1589 271
rect 1635 225 1713 271
rect 1759 225 1837 271
rect 1883 225 1961 271
rect 2007 225 2085 271
rect 2131 225 2209 271
rect 2255 225 2333 271
rect 2379 225 2457 271
rect 2503 225 2581 271
rect 2627 225 2705 271
rect 2751 225 2829 271
rect 2875 225 2953 271
rect 2999 225 3077 271
rect 3123 225 3201 271
rect 3247 225 3325 271
rect 3371 225 3449 271
rect 3495 225 3573 271
rect 3619 225 3697 271
rect 3743 225 3821 271
rect 3867 225 3945 271
rect 3991 225 4069 271
rect 4115 225 4193 271
rect 4239 225 4317 271
rect 4363 225 4441 271
rect 4487 225 4565 271
rect 4611 225 4689 271
rect 4735 225 4813 271
rect 4859 225 4937 271
rect 4983 225 5061 271
rect 5107 225 5185 271
rect 5231 225 5309 271
rect 5355 225 5433 271
rect 5479 225 5557 271
rect 5603 225 5681 271
rect 5727 225 5805 271
rect 5851 225 5929 271
rect 5975 225 6053 271
rect 6099 225 6177 271
rect 6223 225 6301 271
rect 6347 225 6425 271
rect 6471 225 6549 271
rect 6595 225 6673 271
rect 6719 225 6797 271
rect 6843 225 6921 271
rect 6967 225 7045 271
rect 7091 225 7169 271
rect 7215 225 7293 271
rect 7339 225 7417 271
rect 7463 225 7541 271
rect 7587 225 7665 271
rect 7711 225 7789 271
rect 7835 225 7913 271
rect 7959 225 8037 271
rect 8083 225 8161 271
rect 8207 225 8285 271
rect 8331 225 8409 271
rect 8455 225 8533 271
rect 8579 225 8657 271
rect 8703 225 8781 271
rect 8827 225 8905 271
rect 8951 225 9029 271
rect 9075 225 9153 271
rect 9199 225 9277 271
rect 9323 225 9401 271
rect 9447 225 9525 271
rect 9571 225 9649 271
rect 9695 225 9773 271
rect 9819 225 9897 271
rect 9943 225 10021 271
rect 10067 225 10145 271
rect 10191 225 10269 271
rect 10315 225 10393 271
rect 10439 225 10517 271
rect 10563 225 10641 271
rect 10687 225 10765 271
rect 10811 225 10889 271
rect 10935 225 11013 271
rect 11059 225 11137 271
rect 11183 225 11261 271
rect 11307 225 11385 271
rect 11431 225 11509 271
rect 11555 225 11633 271
rect 11679 225 11757 271
rect 11803 225 11881 271
rect 11927 225 12005 271
rect 12051 225 12129 271
rect 12175 225 12253 271
rect 12299 225 12377 271
rect 12423 225 12501 271
rect 12547 225 12625 271
rect 12671 225 12749 271
rect 12795 225 12873 271
rect 12919 225 12997 271
rect 13043 225 13121 271
rect 13167 225 13245 271
rect 13291 225 13369 271
rect 13415 225 13493 271
rect 13539 225 13617 271
rect 13663 225 13741 271
rect 13787 225 13865 271
rect 13911 225 13989 271
rect 14035 225 14113 271
rect 14159 225 14237 271
rect 14283 225 14361 271
rect 14407 225 14485 271
rect 14531 225 14609 271
rect 14655 225 14733 271
rect 14779 225 14857 271
rect 14903 225 14981 271
rect 15027 225 15105 271
rect 15151 225 15229 271
rect 15275 225 15353 271
rect 15399 225 15477 271
rect 15523 225 15601 271
rect 15647 225 15725 271
rect 15771 225 15849 271
rect 15895 225 15973 271
rect 16019 225 16097 271
rect 16143 225 16221 271
rect 16267 225 16345 271
rect 16391 225 16469 271
rect 16515 225 16593 271
rect 16639 225 16717 271
rect 16763 225 16841 271
rect 16887 225 16965 271
rect 17011 225 17089 271
rect 17135 225 17213 271
rect 17259 225 17337 271
rect 17383 225 17461 271
rect 17507 225 17585 271
rect 17631 225 17709 271
rect 17755 225 17833 271
rect 17879 225 17957 271
rect 18003 225 18081 271
rect 18127 225 18205 271
rect 18251 225 18329 271
rect 18375 225 18453 271
rect 18499 225 18577 271
rect 18623 225 18701 271
rect 18747 225 18825 271
rect 18871 225 18949 271
rect 18995 225 19073 271
rect 19119 225 19197 271
rect 19243 225 19321 271
rect 19367 225 19445 271
rect 19491 225 19569 271
rect 19615 225 19693 271
rect 19739 225 19817 271
rect 19863 225 19941 271
rect 19987 225 20065 271
rect 20111 225 20189 271
rect 20235 225 20313 271
rect 20359 225 20437 271
rect 20483 225 20561 271
rect 20607 225 20685 271
rect 20731 225 20809 271
rect 20855 225 20933 271
rect 20979 225 21057 271
rect 21103 225 21181 271
rect 21227 225 21305 271
rect 21351 225 21429 271
rect 21475 225 21553 271
rect 21599 225 21677 271
rect 21723 225 21801 271
rect 21847 225 21925 271
rect 21971 225 22049 271
rect 22095 225 22173 271
rect 22219 225 22297 271
rect 22343 225 22421 271
rect 22467 225 22545 271
rect 22591 225 22669 271
rect 22715 225 22793 271
rect 22839 225 22917 271
rect 22963 225 23041 271
rect 23087 225 23165 271
rect 23211 225 23289 271
rect 23335 225 23413 271
rect 23459 225 23537 271
rect 23583 225 23661 271
rect 23707 225 23785 271
rect 23831 225 23909 271
rect 23955 225 24033 271
rect 24079 225 24157 271
rect 24203 225 24281 271
rect 24327 225 24405 271
rect 24451 225 24529 271
rect 24575 225 24653 271
rect 24699 225 24777 271
rect 24823 225 24901 271
rect 24947 225 25025 271
rect 25071 225 25149 271
rect 25195 225 25273 271
rect 25319 225 25397 271
rect 25443 225 25521 271
rect 25567 225 25645 271
rect 25691 225 25769 271
rect 25815 225 25893 271
rect 25939 225 26017 271
rect 26063 225 26141 271
rect 26187 225 26265 271
rect 26311 225 26389 271
rect 26435 225 26513 271
rect 26559 225 26637 271
rect 26683 225 26761 271
rect 26807 225 26885 271
rect 26931 225 27009 271
rect 27055 225 27133 271
rect 27179 225 27257 271
rect 27303 225 27381 271
rect 27427 225 27505 271
rect 27551 225 27629 271
rect 27675 225 27753 271
rect 27799 225 27877 271
rect 27923 225 28001 271
rect 28047 225 28125 271
rect 28171 225 28249 271
rect 28295 225 28373 271
rect 28419 225 28497 271
rect 28543 225 28621 271
rect 28667 225 28745 271
rect 28791 225 28869 271
rect 28915 225 28993 271
rect 29039 225 29117 271
rect 29163 225 29241 271
rect 29287 225 29365 271
rect 29411 225 29489 271
rect 29535 225 29613 271
rect 29659 225 29737 271
rect 29783 225 29861 271
rect 29907 225 29985 271
rect 30031 225 30109 271
rect 30155 225 30233 271
rect 30279 225 30357 271
rect 30403 225 30481 271
rect 30527 225 30605 271
rect 30651 225 30729 271
rect 30775 225 30853 271
rect 30899 225 30977 271
rect 31023 225 31101 271
rect 31147 225 31225 271
rect 31271 225 31349 271
rect 31395 225 31473 271
rect 31519 225 31597 271
rect 31643 225 31721 271
rect 31767 225 31845 271
rect 31891 225 31969 271
rect 32015 225 32093 271
rect 32139 225 32217 271
rect 32263 225 32341 271
rect 32387 225 32465 271
rect 32511 225 32589 271
rect 32635 225 32713 271
rect 32759 225 32837 271
rect 32883 225 32961 271
rect 33007 225 33085 271
rect 33131 225 33209 271
rect 33255 225 33333 271
rect 33379 225 33457 271
rect 33503 225 33581 271
rect 33627 225 33705 271
rect 33751 225 33829 271
rect 33875 225 33953 271
rect 33999 225 34077 271
rect 34123 225 34201 271
rect 34247 225 34325 271
rect 34371 225 34449 271
rect 34495 225 34573 271
rect 34619 225 34697 271
rect 34743 225 34821 271
rect 34867 225 34945 271
rect 34991 225 35069 271
rect 35115 225 35193 271
rect 35239 225 35317 271
rect 35363 225 35441 271
rect 35487 225 35565 271
rect 35611 225 35689 271
rect 35735 225 35813 271
rect 35859 225 35937 271
rect 35983 225 36061 271
rect 36107 225 36185 271
rect 36231 225 36309 271
rect 36355 225 36433 271
rect 36479 225 36557 271
rect 36603 225 36681 271
rect 36727 225 36805 271
rect 36851 225 36929 271
rect 36975 225 37053 271
rect 37099 225 37177 271
rect 37223 225 37301 271
rect 37347 225 37425 271
rect 37471 225 37549 271
rect 37595 225 37673 271
rect 37719 225 37797 271
rect 37843 225 37921 271
rect 37967 225 38045 271
rect 38091 225 38169 271
rect 38215 225 38293 271
rect 38339 225 38417 271
rect 38463 225 38541 271
rect 38587 225 38665 271
rect 38711 225 38789 271
rect 38835 225 38913 271
rect 38959 225 39037 271
rect 39083 225 39161 271
rect 39207 225 39285 271
rect 39331 225 39409 271
rect 39455 225 39533 271
rect 39579 225 39657 271
rect 39703 225 39781 271
rect 39827 225 39905 271
rect 39951 225 40029 271
rect 40075 225 40153 271
rect 40199 225 40277 271
rect 40323 225 40401 271
rect 40447 225 40525 271
rect 40571 225 40649 271
rect 40695 225 40773 271
rect 40819 225 40897 271
rect 40943 225 41021 271
rect 41067 225 41145 271
rect 41191 225 41269 271
rect 41315 225 41393 271
rect 41439 225 41517 271
rect 41563 225 41641 271
rect 41687 225 41765 271
rect 41811 225 41889 271
rect 41935 225 42013 271
rect 42059 225 42137 271
rect 42183 225 42261 271
rect 42307 225 42385 271
rect 42431 225 42509 271
rect 42555 225 42633 271
rect 42679 225 42757 271
rect 42803 225 42881 271
rect 42927 225 43005 271
rect 43051 225 43129 271
rect 43175 225 43253 271
rect 43299 225 43377 271
rect 43423 225 43501 271
rect 43547 225 43625 271
rect 43671 225 43749 271
rect 43795 225 43873 271
rect 43919 225 43997 271
rect 44043 225 44121 271
rect 44167 225 44245 271
rect 44291 225 44369 271
rect 44415 225 44493 271
rect 44539 225 44617 271
rect 44663 225 44741 271
rect 44787 225 44865 271
rect 44911 225 44989 271
rect 45035 225 45113 271
rect 45159 225 45237 271
rect 45283 225 45361 271
rect 45407 225 45485 271
rect 45531 225 45609 271
rect 45655 225 45733 271
rect 45779 225 45857 271
rect 45903 225 45981 271
rect 46027 225 46105 271
rect 46151 225 46229 271
rect 46275 225 46353 271
rect 46399 225 46477 271
rect 46523 225 46601 271
rect 46647 225 46725 271
rect 46771 225 46849 271
rect 46895 225 46973 271
rect 47019 225 47097 271
rect 47143 225 47221 271
rect 47267 225 47345 271
rect 47391 225 47469 271
rect 47515 225 47593 271
rect 47639 225 47717 271
rect 47763 225 47841 271
rect 47887 225 47965 271
rect 48011 225 48089 271
rect 48135 225 48213 271
rect 48259 225 48337 271
rect 48383 225 48461 271
rect 48507 225 48585 271
rect 48631 225 48709 271
rect 48755 225 48833 271
rect 48879 225 48957 271
rect 49003 225 49081 271
rect 49127 225 49205 271
rect 49251 225 49329 271
rect 49375 225 49453 271
rect 49499 225 49577 271
rect 49623 225 49701 271
rect 49747 225 49825 271
rect 49871 225 49949 271
rect 49995 225 50073 271
rect 50119 225 50197 271
rect 50243 225 50321 271
rect 50367 225 50445 271
rect 50491 225 50569 271
rect 50615 225 50693 271
rect 50739 225 50817 271
rect 50863 225 50941 271
rect 50987 225 51065 271
rect 51111 225 51189 271
rect 51235 225 51313 271
rect 51359 225 51437 271
rect 51483 225 51561 271
rect 51607 225 51685 271
rect 51731 225 51809 271
rect 51855 225 51933 271
rect 51979 225 52057 271
rect 52103 225 52181 271
rect 52227 225 52305 271
rect 52351 225 52429 271
rect 52475 225 52553 271
rect 52599 225 52677 271
rect 52723 225 52801 271
rect 52847 225 52925 271
rect 52971 225 53049 271
rect 53095 225 53173 271
rect 53219 225 53297 271
rect 53343 225 53421 271
rect 53467 225 53545 271
rect 53591 225 53669 271
rect 53715 225 53793 271
rect 53839 225 53917 271
rect 53963 225 54041 271
rect 54087 225 54165 271
rect 54211 225 54289 271
rect 54335 225 54413 271
rect 54459 225 54537 271
rect 54583 225 54661 271
rect 54707 225 54785 271
rect 54831 225 54909 271
rect 54955 225 55033 271
rect 55079 225 55157 271
rect 55203 225 55281 271
rect 55327 225 55405 271
rect 55451 225 55529 271
rect 55575 225 55653 271
rect 55699 225 55777 271
rect 55823 225 55901 271
rect 55947 225 56025 271
rect 56071 225 56149 271
rect 56195 225 56273 271
rect 56319 225 56397 271
rect 56443 225 56521 271
rect 56567 225 56645 271
rect 56691 225 56769 271
rect 56815 225 56893 271
rect 56939 225 57017 271
rect 57063 225 57141 271
rect 57187 225 57265 271
rect 57311 225 57389 271
rect 57435 225 57513 271
rect 57559 225 57637 271
rect 57683 225 57761 271
rect 57807 225 57885 271
rect 57931 225 58009 271
rect 58055 225 58133 271
rect 58179 225 58257 271
rect 58303 225 58381 271
rect 58427 225 58505 271
rect 58551 225 58629 271
rect 58675 225 58753 271
rect 58799 225 58877 271
rect 58923 225 59001 271
rect 59047 225 59125 271
rect 59171 225 59249 271
rect 59295 225 59373 271
rect 59419 225 59497 271
rect 59543 225 59621 271
rect 59667 225 59745 271
rect 59791 225 59869 271
rect 59915 225 59993 271
rect 60039 225 60117 271
rect 60163 225 60241 271
rect 60287 225 60365 271
rect 60411 225 60489 271
rect 60535 225 60613 271
rect 60659 225 60737 271
rect 60783 225 60861 271
rect 60907 225 60985 271
rect 61031 225 61109 271
rect 61155 225 61233 271
rect 61279 225 61357 271
rect 61403 225 61481 271
rect 61527 225 61605 271
rect 61651 225 61729 271
rect 61775 225 61853 271
rect 61899 225 61977 271
rect 62023 225 62101 271
rect 62147 225 62225 271
rect 62271 225 62349 271
rect 62395 225 62473 271
rect 62519 225 62597 271
rect 62643 225 62721 271
rect 62767 225 62845 271
rect 62891 225 62969 271
rect 63015 225 63093 271
rect 63139 225 63217 271
rect 63263 225 63341 271
rect 63387 225 63465 271
rect 63511 225 63589 271
rect 63635 225 63713 271
rect 63759 225 63837 271
rect 63883 225 63961 271
rect 64007 225 64085 271
rect 64131 225 64209 271
rect 64255 225 64333 271
rect 64379 225 64457 271
rect 64503 225 64581 271
rect 64627 225 64705 271
rect 64751 225 64829 271
rect 64875 225 64953 271
rect 64999 225 65077 271
rect 65123 225 65201 271
rect 65247 225 65325 271
rect 65371 225 65449 271
rect 65495 225 65573 271
rect 65619 225 65697 271
rect 65743 225 65821 271
rect 65867 225 65945 271
rect 65991 225 66069 271
rect 66115 225 66193 271
rect 66239 225 66317 271
rect 66363 225 66441 271
rect 66487 225 66565 271
rect 66611 225 66689 271
rect 66735 225 66813 271
rect 66859 225 66937 271
rect 66983 225 67061 271
rect 67107 225 67185 271
rect 67231 225 67309 271
rect 67355 225 67433 271
rect 67479 225 67557 271
rect 67603 225 67681 271
rect 67727 225 67805 271
rect 67851 225 67929 271
rect 67975 225 68053 271
rect 68099 225 68177 271
rect 68223 225 68301 271
rect 68347 225 68425 271
rect 68471 225 68549 271
rect 68595 225 68673 271
rect 68719 225 68797 271
rect 68843 225 68921 271
rect 68967 225 69045 271
rect 69091 225 69169 271
rect 69215 225 69293 271
rect 69339 225 69417 271
rect 69463 225 69541 271
rect 69587 225 69665 271
rect 69711 225 69789 271
rect 69835 225 69913 271
rect 69959 225 70037 271
rect 70083 225 70161 271
rect 70207 225 70285 271
rect 70331 225 70409 271
rect 70455 225 70533 271
rect 70579 225 70657 271
rect 70703 225 70781 271
rect 70827 225 70905 271
rect 70951 225 71029 271
rect 71075 225 71153 271
rect 71199 225 71277 271
rect 71323 225 71401 271
rect 71447 225 71525 271
rect 71571 225 71649 271
rect 71695 225 71773 271
rect 71819 225 71897 271
rect 71943 225 72021 271
rect 72067 225 72145 271
rect 72191 225 72269 271
rect 72315 225 72393 271
rect 72439 225 72517 271
rect 72563 225 72641 271
rect 72687 225 72765 271
rect 72811 225 72889 271
rect 72935 225 73013 271
rect 73059 225 73137 271
rect 73183 225 73261 271
rect 73307 225 73385 271
rect 73431 225 73509 271
rect 73555 225 73633 271
rect 73679 225 73757 271
rect 73803 225 73881 271
rect 73927 225 74005 271
rect 74051 225 74129 271
rect 74175 225 74253 271
rect 74299 225 74377 271
rect 74423 225 74501 271
rect 74547 225 74625 271
rect 74671 225 74749 271
rect 74795 225 74873 271
rect 74919 225 74997 271
rect 75043 225 75121 271
rect 75167 225 75245 271
rect 75291 225 75369 271
rect 75415 225 75493 271
rect 75539 225 75617 271
rect 75663 225 75741 271
rect 75787 225 75865 271
rect 75911 225 75989 271
rect 76035 225 76113 271
rect 76159 225 76237 271
rect 76283 225 76361 271
rect 76407 225 76485 271
rect 76531 225 76609 271
rect 76655 225 76733 271
rect 76779 225 76857 271
rect 76903 225 76981 271
rect 77027 225 77105 271
rect 77151 225 77229 271
rect 77275 225 77353 271
rect 77399 225 77477 271
rect 77523 225 77601 271
rect 77647 225 77725 271
rect 77771 225 77849 271
rect 77895 225 77973 271
rect 78019 225 78097 271
rect 78143 225 78221 271
rect 78267 225 78345 271
rect 78391 225 78469 271
rect 78515 225 78593 271
rect 78639 225 78717 271
rect 78763 225 78841 271
rect 78887 225 78965 271
rect 79011 225 79089 271
rect 79135 225 79213 271
rect 79259 225 79337 271
rect 79383 225 79461 271
rect 79507 225 79585 271
rect 79631 225 79709 271
rect 79755 225 79833 271
rect 79879 225 79957 271
rect 80003 225 80081 271
rect 80127 225 80205 271
rect 80251 225 80329 271
rect 80375 225 80453 271
rect 80499 225 80577 271
rect 80623 225 80701 271
rect 80747 225 80825 271
rect 80871 225 80949 271
rect 80995 225 81073 271
rect 81119 225 81197 271
rect 81243 225 81321 271
rect 81367 225 81445 271
rect 81491 225 81569 271
rect 81615 225 81693 271
rect 81739 225 81817 271
rect 81863 225 81941 271
rect 81987 225 82065 271
rect 82111 225 82189 271
rect 82235 225 82313 271
rect 82359 225 82437 271
rect 82483 225 82561 271
rect 82607 225 82685 271
rect 82731 225 82809 271
rect 82855 225 82933 271
rect 82979 225 83057 271
rect 83103 225 83181 271
rect 83227 225 83305 271
rect 83351 225 83429 271
rect 83475 225 83553 271
rect 83599 225 83677 271
rect 83723 225 83801 271
rect 83847 225 83925 271
rect 83971 225 84049 271
rect 84095 225 84173 271
rect 84219 225 84297 271
rect 84343 225 84421 271
rect 84467 225 84545 271
rect 84591 225 84669 271
rect 84715 225 84793 271
rect 84839 225 84917 271
rect 84963 225 85041 271
rect 85087 225 85165 271
rect 85211 225 85289 271
rect 85335 225 85413 271
rect 85459 225 85537 271
rect 85583 225 85602 271
rect -42 147 85602 225
rect -42 101 -23 147
rect 23 101 101 147
rect 147 101 225 147
rect 271 101 349 147
rect 395 101 473 147
rect 519 101 597 147
rect 643 101 721 147
rect 767 101 845 147
rect 891 101 969 147
rect 1015 101 1093 147
rect 1139 101 1217 147
rect 1263 101 1341 147
rect 1387 101 1465 147
rect 1511 101 1589 147
rect 1635 101 1713 147
rect 1759 101 1837 147
rect 1883 101 1961 147
rect 2007 101 2085 147
rect 2131 101 2209 147
rect 2255 101 2333 147
rect 2379 101 2457 147
rect 2503 101 2581 147
rect 2627 101 2705 147
rect 2751 101 2829 147
rect 2875 101 2953 147
rect 2999 101 3077 147
rect 3123 101 3201 147
rect 3247 101 3325 147
rect 3371 101 3449 147
rect 3495 101 3573 147
rect 3619 101 3697 147
rect 3743 101 3821 147
rect 3867 101 3945 147
rect 3991 101 4069 147
rect 4115 101 4193 147
rect 4239 101 4317 147
rect 4363 101 4441 147
rect 4487 101 4565 147
rect 4611 101 4689 147
rect 4735 101 4813 147
rect 4859 101 4937 147
rect 4983 101 5061 147
rect 5107 101 5185 147
rect 5231 101 5309 147
rect 5355 101 5433 147
rect 5479 101 5557 147
rect 5603 101 5681 147
rect 5727 101 5805 147
rect 5851 101 5929 147
rect 5975 101 6053 147
rect 6099 101 6177 147
rect 6223 101 6301 147
rect 6347 101 6425 147
rect 6471 101 6549 147
rect 6595 101 6673 147
rect 6719 101 6797 147
rect 6843 101 6921 147
rect 6967 101 7045 147
rect 7091 101 7169 147
rect 7215 101 7293 147
rect 7339 101 7417 147
rect 7463 101 7541 147
rect 7587 101 7665 147
rect 7711 101 7789 147
rect 7835 101 7913 147
rect 7959 101 8037 147
rect 8083 101 8161 147
rect 8207 101 8285 147
rect 8331 101 8409 147
rect 8455 101 8533 147
rect 8579 101 8657 147
rect 8703 101 8781 147
rect 8827 101 8905 147
rect 8951 101 9029 147
rect 9075 101 9153 147
rect 9199 101 9277 147
rect 9323 101 9401 147
rect 9447 101 9525 147
rect 9571 101 9649 147
rect 9695 101 9773 147
rect 9819 101 9897 147
rect 9943 101 10021 147
rect 10067 101 10145 147
rect 10191 101 10269 147
rect 10315 101 10393 147
rect 10439 101 10517 147
rect 10563 101 10641 147
rect 10687 101 10765 147
rect 10811 101 10889 147
rect 10935 101 11013 147
rect 11059 101 11137 147
rect 11183 101 11261 147
rect 11307 101 11385 147
rect 11431 101 11509 147
rect 11555 101 11633 147
rect 11679 101 11757 147
rect 11803 101 11881 147
rect 11927 101 12005 147
rect 12051 101 12129 147
rect 12175 101 12253 147
rect 12299 101 12377 147
rect 12423 101 12501 147
rect 12547 101 12625 147
rect 12671 101 12749 147
rect 12795 101 12873 147
rect 12919 101 12997 147
rect 13043 101 13121 147
rect 13167 101 13245 147
rect 13291 101 13369 147
rect 13415 101 13493 147
rect 13539 101 13617 147
rect 13663 101 13741 147
rect 13787 101 13865 147
rect 13911 101 13989 147
rect 14035 101 14113 147
rect 14159 101 14237 147
rect 14283 101 14361 147
rect 14407 101 14485 147
rect 14531 101 14609 147
rect 14655 101 14733 147
rect 14779 101 14857 147
rect 14903 101 14981 147
rect 15027 101 15105 147
rect 15151 101 15229 147
rect 15275 101 15353 147
rect 15399 101 15477 147
rect 15523 101 15601 147
rect 15647 101 15725 147
rect 15771 101 15849 147
rect 15895 101 15973 147
rect 16019 101 16097 147
rect 16143 101 16221 147
rect 16267 101 16345 147
rect 16391 101 16469 147
rect 16515 101 16593 147
rect 16639 101 16717 147
rect 16763 101 16841 147
rect 16887 101 16965 147
rect 17011 101 17089 147
rect 17135 101 17213 147
rect 17259 101 17337 147
rect 17383 101 17461 147
rect 17507 101 17585 147
rect 17631 101 17709 147
rect 17755 101 17833 147
rect 17879 101 17957 147
rect 18003 101 18081 147
rect 18127 101 18205 147
rect 18251 101 18329 147
rect 18375 101 18453 147
rect 18499 101 18577 147
rect 18623 101 18701 147
rect 18747 101 18825 147
rect 18871 101 18949 147
rect 18995 101 19073 147
rect 19119 101 19197 147
rect 19243 101 19321 147
rect 19367 101 19445 147
rect 19491 101 19569 147
rect 19615 101 19693 147
rect 19739 101 19817 147
rect 19863 101 19941 147
rect 19987 101 20065 147
rect 20111 101 20189 147
rect 20235 101 20313 147
rect 20359 101 20437 147
rect 20483 101 20561 147
rect 20607 101 20685 147
rect 20731 101 20809 147
rect 20855 101 20933 147
rect 20979 101 21057 147
rect 21103 101 21181 147
rect 21227 101 21305 147
rect 21351 101 21429 147
rect 21475 101 21553 147
rect 21599 101 21677 147
rect 21723 101 21801 147
rect 21847 101 21925 147
rect 21971 101 22049 147
rect 22095 101 22173 147
rect 22219 101 22297 147
rect 22343 101 22421 147
rect 22467 101 22545 147
rect 22591 101 22669 147
rect 22715 101 22793 147
rect 22839 101 22917 147
rect 22963 101 23041 147
rect 23087 101 23165 147
rect 23211 101 23289 147
rect 23335 101 23413 147
rect 23459 101 23537 147
rect 23583 101 23661 147
rect 23707 101 23785 147
rect 23831 101 23909 147
rect 23955 101 24033 147
rect 24079 101 24157 147
rect 24203 101 24281 147
rect 24327 101 24405 147
rect 24451 101 24529 147
rect 24575 101 24653 147
rect 24699 101 24777 147
rect 24823 101 24901 147
rect 24947 101 25025 147
rect 25071 101 25149 147
rect 25195 101 25273 147
rect 25319 101 25397 147
rect 25443 101 25521 147
rect 25567 101 25645 147
rect 25691 101 25769 147
rect 25815 101 25893 147
rect 25939 101 26017 147
rect 26063 101 26141 147
rect 26187 101 26265 147
rect 26311 101 26389 147
rect 26435 101 26513 147
rect 26559 101 26637 147
rect 26683 101 26761 147
rect 26807 101 26885 147
rect 26931 101 27009 147
rect 27055 101 27133 147
rect 27179 101 27257 147
rect 27303 101 27381 147
rect 27427 101 27505 147
rect 27551 101 27629 147
rect 27675 101 27753 147
rect 27799 101 27877 147
rect 27923 101 28001 147
rect 28047 101 28125 147
rect 28171 101 28249 147
rect 28295 101 28373 147
rect 28419 101 28497 147
rect 28543 101 28621 147
rect 28667 101 28745 147
rect 28791 101 28869 147
rect 28915 101 28993 147
rect 29039 101 29117 147
rect 29163 101 29241 147
rect 29287 101 29365 147
rect 29411 101 29489 147
rect 29535 101 29613 147
rect 29659 101 29737 147
rect 29783 101 29861 147
rect 29907 101 29985 147
rect 30031 101 30109 147
rect 30155 101 30233 147
rect 30279 101 30357 147
rect 30403 101 30481 147
rect 30527 101 30605 147
rect 30651 101 30729 147
rect 30775 101 30853 147
rect 30899 101 30977 147
rect 31023 101 31101 147
rect 31147 101 31225 147
rect 31271 101 31349 147
rect 31395 101 31473 147
rect 31519 101 31597 147
rect 31643 101 31721 147
rect 31767 101 31845 147
rect 31891 101 31969 147
rect 32015 101 32093 147
rect 32139 101 32217 147
rect 32263 101 32341 147
rect 32387 101 32465 147
rect 32511 101 32589 147
rect 32635 101 32713 147
rect 32759 101 32837 147
rect 32883 101 32961 147
rect 33007 101 33085 147
rect 33131 101 33209 147
rect 33255 101 33333 147
rect 33379 101 33457 147
rect 33503 101 33581 147
rect 33627 101 33705 147
rect 33751 101 33829 147
rect 33875 101 33953 147
rect 33999 101 34077 147
rect 34123 101 34201 147
rect 34247 101 34325 147
rect 34371 101 34449 147
rect 34495 101 34573 147
rect 34619 101 34697 147
rect 34743 101 34821 147
rect 34867 101 34945 147
rect 34991 101 35069 147
rect 35115 101 35193 147
rect 35239 101 35317 147
rect 35363 101 35441 147
rect 35487 101 35565 147
rect 35611 101 35689 147
rect 35735 101 35813 147
rect 35859 101 35937 147
rect 35983 101 36061 147
rect 36107 101 36185 147
rect 36231 101 36309 147
rect 36355 101 36433 147
rect 36479 101 36557 147
rect 36603 101 36681 147
rect 36727 101 36805 147
rect 36851 101 36929 147
rect 36975 101 37053 147
rect 37099 101 37177 147
rect 37223 101 37301 147
rect 37347 101 37425 147
rect 37471 101 37549 147
rect 37595 101 37673 147
rect 37719 101 37797 147
rect 37843 101 37921 147
rect 37967 101 38045 147
rect 38091 101 38169 147
rect 38215 101 38293 147
rect 38339 101 38417 147
rect 38463 101 38541 147
rect 38587 101 38665 147
rect 38711 101 38789 147
rect 38835 101 38913 147
rect 38959 101 39037 147
rect 39083 101 39161 147
rect 39207 101 39285 147
rect 39331 101 39409 147
rect 39455 101 39533 147
rect 39579 101 39657 147
rect 39703 101 39781 147
rect 39827 101 39905 147
rect 39951 101 40029 147
rect 40075 101 40153 147
rect 40199 101 40277 147
rect 40323 101 40401 147
rect 40447 101 40525 147
rect 40571 101 40649 147
rect 40695 101 40773 147
rect 40819 101 40897 147
rect 40943 101 41021 147
rect 41067 101 41145 147
rect 41191 101 41269 147
rect 41315 101 41393 147
rect 41439 101 41517 147
rect 41563 101 41641 147
rect 41687 101 41765 147
rect 41811 101 41889 147
rect 41935 101 42013 147
rect 42059 101 42137 147
rect 42183 101 42261 147
rect 42307 101 42385 147
rect 42431 101 42509 147
rect 42555 101 42633 147
rect 42679 101 42757 147
rect 42803 101 42881 147
rect 42927 101 43005 147
rect 43051 101 43129 147
rect 43175 101 43253 147
rect 43299 101 43377 147
rect 43423 101 43501 147
rect 43547 101 43625 147
rect 43671 101 43749 147
rect 43795 101 43873 147
rect 43919 101 43997 147
rect 44043 101 44121 147
rect 44167 101 44245 147
rect 44291 101 44369 147
rect 44415 101 44493 147
rect 44539 101 44617 147
rect 44663 101 44741 147
rect 44787 101 44865 147
rect 44911 101 44989 147
rect 45035 101 45113 147
rect 45159 101 45237 147
rect 45283 101 45361 147
rect 45407 101 45485 147
rect 45531 101 45609 147
rect 45655 101 45733 147
rect 45779 101 45857 147
rect 45903 101 45981 147
rect 46027 101 46105 147
rect 46151 101 46229 147
rect 46275 101 46353 147
rect 46399 101 46477 147
rect 46523 101 46601 147
rect 46647 101 46725 147
rect 46771 101 46849 147
rect 46895 101 46973 147
rect 47019 101 47097 147
rect 47143 101 47221 147
rect 47267 101 47345 147
rect 47391 101 47469 147
rect 47515 101 47593 147
rect 47639 101 47717 147
rect 47763 101 47841 147
rect 47887 101 47965 147
rect 48011 101 48089 147
rect 48135 101 48213 147
rect 48259 101 48337 147
rect 48383 101 48461 147
rect 48507 101 48585 147
rect 48631 101 48709 147
rect 48755 101 48833 147
rect 48879 101 48957 147
rect 49003 101 49081 147
rect 49127 101 49205 147
rect 49251 101 49329 147
rect 49375 101 49453 147
rect 49499 101 49577 147
rect 49623 101 49701 147
rect 49747 101 49825 147
rect 49871 101 49949 147
rect 49995 101 50073 147
rect 50119 101 50197 147
rect 50243 101 50321 147
rect 50367 101 50445 147
rect 50491 101 50569 147
rect 50615 101 50693 147
rect 50739 101 50817 147
rect 50863 101 50941 147
rect 50987 101 51065 147
rect 51111 101 51189 147
rect 51235 101 51313 147
rect 51359 101 51437 147
rect 51483 101 51561 147
rect 51607 101 51685 147
rect 51731 101 51809 147
rect 51855 101 51933 147
rect 51979 101 52057 147
rect 52103 101 52181 147
rect 52227 101 52305 147
rect 52351 101 52429 147
rect 52475 101 52553 147
rect 52599 101 52677 147
rect 52723 101 52801 147
rect 52847 101 52925 147
rect 52971 101 53049 147
rect 53095 101 53173 147
rect 53219 101 53297 147
rect 53343 101 53421 147
rect 53467 101 53545 147
rect 53591 101 53669 147
rect 53715 101 53793 147
rect 53839 101 53917 147
rect 53963 101 54041 147
rect 54087 101 54165 147
rect 54211 101 54289 147
rect 54335 101 54413 147
rect 54459 101 54537 147
rect 54583 101 54661 147
rect 54707 101 54785 147
rect 54831 101 54909 147
rect 54955 101 55033 147
rect 55079 101 55157 147
rect 55203 101 55281 147
rect 55327 101 55405 147
rect 55451 101 55529 147
rect 55575 101 55653 147
rect 55699 101 55777 147
rect 55823 101 55901 147
rect 55947 101 56025 147
rect 56071 101 56149 147
rect 56195 101 56273 147
rect 56319 101 56397 147
rect 56443 101 56521 147
rect 56567 101 56645 147
rect 56691 101 56769 147
rect 56815 101 56893 147
rect 56939 101 57017 147
rect 57063 101 57141 147
rect 57187 101 57265 147
rect 57311 101 57389 147
rect 57435 101 57513 147
rect 57559 101 57637 147
rect 57683 101 57761 147
rect 57807 101 57885 147
rect 57931 101 58009 147
rect 58055 101 58133 147
rect 58179 101 58257 147
rect 58303 101 58381 147
rect 58427 101 58505 147
rect 58551 101 58629 147
rect 58675 101 58753 147
rect 58799 101 58877 147
rect 58923 101 59001 147
rect 59047 101 59125 147
rect 59171 101 59249 147
rect 59295 101 59373 147
rect 59419 101 59497 147
rect 59543 101 59621 147
rect 59667 101 59745 147
rect 59791 101 59869 147
rect 59915 101 59993 147
rect 60039 101 60117 147
rect 60163 101 60241 147
rect 60287 101 60365 147
rect 60411 101 60489 147
rect 60535 101 60613 147
rect 60659 101 60737 147
rect 60783 101 60861 147
rect 60907 101 60985 147
rect 61031 101 61109 147
rect 61155 101 61233 147
rect 61279 101 61357 147
rect 61403 101 61481 147
rect 61527 101 61605 147
rect 61651 101 61729 147
rect 61775 101 61853 147
rect 61899 101 61977 147
rect 62023 101 62101 147
rect 62147 101 62225 147
rect 62271 101 62349 147
rect 62395 101 62473 147
rect 62519 101 62597 147
rect 62643 101 62721 147
rect 62767 101 62845 147
rect 62891 101 62969 147
rect 63015 101 63093 147
rect 63139 101 63217 147
rect 63263 101 63341 147
rect 63387 101 63465 147
rect 63511 101 63589 147
rect 63635 101 63713 147
rect 63759 101 63837 147
rect 63883 101 63961 147
rect 64007 101 64085 147
rect 64131 101 64209 147
rect 64255 101 64333 147
rect 64379 101 64457 147
rect 64503 101 64581 147
rect 64627 101 64705 147
rect 64751 101 64829 147
rect 64875 101 64953 147
rect 64999 101 65077 147
rect 65123 101 65201 147
rect 65247 101 65325 147
rect 65371 101 65449 147
rect 65495 101 65573 147
rect 65619 101 65697 147
rect 65743 101 65821 147
rect 65867 101 65945 147
rect 65991 101 66069 147
rect 66115 101 66193 147
rect 66239 101 66317 147
rect 66363 101 66441 147
rect 66487 101 66565 147
rect 66611 101 66689 147
rect 66735 101 66813 147
rect 66859 101 66937 147
rect 66983 101 67061 147
rect 67107 101 67185 147
rect 67231 101 67309 147
rect 67355 101 67433 147
rect 67479 101 67557 147
rect 67603 101 67681 147
rect 67727 101 67805 147
rect 67851 101 67929 147
rect 67975 101 68053 147
rect 68099 101 68177 147
rect 68223 101 68301 147
rect 68347 101 68425 147
rect 68471 101 68549 147
rect 68595 101 68673 147
rect 68719 101 68797 147
rect 68843 101 68921 147
rect 68967 101 69045 147
rect 69091 101 69169 147
rect 69215 101 69293 147
rect 69339 101 69417 147
rect 69463 101 69541 147
rect 69587 101 69665 147
rect 69711 101 69789 147
rect 69835 101 69913 147
rect 69959 101 70037 147
rect 70083 101 70161 147
rect 70207 101 70285 147
rect 70331 101 70409 147
rect 70455 101 70533 147
rect 70579 101 70657 147
rect 70703 101 70781 147
rect 70827 101 70905 147
rect 70951 101 71029 147
rect 71075 101 71153 147
rect 71199 101 71277 147
rect 71323 101 71401 147
rect 71447 101 71525 147
rect 71571 101 71649 147
rect 71695 101 71773 147
rect 71819 101 71897 147
rect 71943 101 72021 147
rect 72067 101 72145 147
rect 72191 101 72269 147
rect 72315 101 72393 147
rect 72439 101 72517 147
rect 72563 101 72641 147
rect 72687 101 72765 147
rect 72811 101 72889 147
rect 72935 101 73013 147
rect 73059 101 73137 147
rect 73183 101 73261 147
rect 73307 101 73385 147
rect 73431 101 73509 147
rect 73555 101 73633 147
rect 73679 101 73757 147
rect 73803 101 73881 147
rect 73927 101 74005 147
rect 74051 101 74129 147
rect 74175 101 74253 147
rect 74299 101 74377 147
rect 74423 101 74501 147
rect 74547 101 74625 147
rect 74671 101 74749 147
rect 74795 101 74873 147
rect 74919 101 74997 147
rect 75043 101 75121 147
rect 75167 101 75245 147
rect 75291 101 75369 147
rect 75415 101 75493 147
rect 75539 101 75617 147
rect 75663 101 75741 147
rect 75787 101 75865 147
rect 75911 101 75989 147
rect 76035 101 76113 147
rect 76159 101 76237 147
rect 76283 101 76361 147
rect 76407 101 76485 147
rect 76531 101 76609 147
rect 76655 101 76733 147
rect 76779 101 76857 147
rect 76903 101 76981 147
rect 77027 101 77105 147
rect 77151 101 77229 147
rect 77275 101 77353 147
rect 77399 101 77477 147
rect 77523 101 77601 147
rect 77647 101 77725 147
rect 77771 101 77849 147
rect 77895 101 77973 147
rect 78019 101 78097 147
rect 78143 101 78221 147
rect 78267 101 78345 147
rect 78391 101 78469 147
rect 78515 101 78593 147
rect 78639 101 78717 147
rect 78763 101 78841 147
rect 78887 101 78965 147
rect 79011 101 79089 147
rect 79135 101 79213 147
rect 79259 101 79337 147
rect 79383 101 79461 147
rect 79507 101 79585 147
rect 79631 101 79709 147
rect 79755 101 79833 147
rect 79879 101 79957 147
rect 80003 101 80081 147
rect 80127 101 80205 147
rect 80251 101 80329 147
rect 80375 101 80453 147
rect 80499 101 80577 147
rect 80623 101 80701 147
rect 80747 101 80825 147
rect 80871 101 80949 147
rect 80995 101 81073 147
rect 81119 101 81197 147
rect 81243 101 81321 147
rect 81367 101 81445 147
rect 81491 101 81569 147
rect 81615 101 81693 147
rect 81739 101 81817 147
rect 81863 101 81941 147
rect 81987 101 82065 147
rect 82111 101 82189 147
rect 82235 101 82313 147
rect 82359 101 82437 147
rect 82483 101 82561 147
rect 82607 101 82685 147
rect 82731 101 82809 147
rect 82855 101 82933 147
rect 82979 101 83057 147
rect 83103 101 83181 147
rect 83227 101 83305 147
rect 83351 101 83429 147
rect 83475 101 83553 147
rect 83599 101 83677 147
rect 83723 101 83801 147
rect 83847 101 83925 147
rect 83971 101 84049 147
rect 84095 101 84173 147
rect 84219 101 84297 147
rect 84343 101 84421 147
rect 84467 101 84545 147
rect 84591 101 84669 147
rect 84715 101 84793 147
rect 84839 101 84917 147
rect 84963 101 85041 147
rect 85087 101 85165 147
rect 85211 101 85289 147
rect 85335 101 85413 147
rect 85459 101 85537 147
rect 85583 101 85602 147
rect -42 23 85602 101
rect -42 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 969 23
rect 1015 -23 1093 23
rect 1139 -23 1217 23
rect 1263 -23 1341 23
rect 1387 -23 1465 23
rect 1511 -23 1589 23
rect 1635 -23 1713 23
rect 1759 -23 1837 23
rect 1883 -23 1961 23
rect 2007 -23 2085 23
rect 2131 -23 2209 23
rect 2255 -23 2333 23
rect 2379 -23 2457 23
rect 2503 -23 2581 23
rect 2627 -23 2705 23
rect 2751 -23 2829 23
rect 2875 -23 2953 23
rect 2999 -23 3077 23
rect 3123 -23 3201 23
rect 3247 -23 3325 23
rect 3371 -23 3449 23
rect 3495 -23 3573 23
rect 3619 -23 3697 23
rect 3743 -23 3821 23
rect 3867 -23 3945 23
rect 3991 -23 4069 23
rect 4115 -23 4193 23
rect 4239 -23 4317 23
rect 4363 -23 4441 23
rect 4487 -23 4565 23
rect 4611 -23 4689 23
rect 4735 -23 4813 23
rect 4859 -23 4937 23
rect 4983 -23 5061 23
rect 5107 -23 5185 23
rect 5231 -23 5309 23
rect 5355 -23 5433 23
rect 5479 -23 5557 23
rect 5603 -23 5681 23
rect 5727 -23 5805 23
rect 5851 -23 5929 23
rect 5975 -23 6053 23
rect 6099 -23 6177 23
rect 6223 -23 6301 23
rect 6347 -23 6425 23
rect 6471 -23 6549 23
rect 6595 -23 6673 23
rect 6719 -23 6797 23
rect 6843 -23 6921 23
rect 6967 -23 7045 23
rect 7091 -23 7169 23
rect 7215 -23 7293 23
rect 7339 -23 7417 23
rect 7463 -23 7541 23
rect 7587 -23 7665 23
rect 7711 -23 7789 23
rect 7835 -23 7913 23
rect 7959 -23 8037 23
rect 8083 -23 8161 23
rect 8207 -23 8285 23
rect 8331 -23 8409 23
rect 8455 -23 8533 23
rect 8579 -23 8657 23
rect 8703 -23 8781 23
rect 8827 -23 8905 23
rect 8951 -23 9029 23
rect 9075 -23 9153 23
rect 9199 -23 9277 23
rect 9323 -23 9401 23
rect 9447 -23 9525 23
rect 9571 -23 9649 23
rect 9695 -23 9773 23
rect 9819 -23 9897 23
rect 9943 -23 10021 23
rect 10067 -23 10145 23
rect 10191 -23 10269 23
rect 10315 -23 10393 23
rect 10439 -23 10517 23
rect 10563 -23 10641 23
rect 10687 -23 10765 23
rect 10811 -23 10889 23
rect 10935 -23 11013 23
rect 11059 -23 11137 23
rect 11183 -23 11261 23
rect 11307 -23 11385 23
rect 11431 -23 11509 23
rect 11555 -23 11633 23
rect 11679 -23 11757 23
rect 11803 -23 11881 23
rect 11927 -23 12005 23
rect 12051 -23 12129 23
rect 12175 -23 12253 23
rect 12299 -23 12377 23
rect 12423 -23 12501 23
rect 12547 -23 12625 23
rect 12671 -23 12749 23
rect 12795 -23 12873 23
rect 12919 -23 12997 23
rect 13043 -23 13121 23
rect 13167 -23 13245 23
rect 13291 -23 13369 23
rect 13415 -23 13493 23
rect 13539 -23 13617 23
rect 13663 -23 13741 23
rect 13787 -23 13865 23
rect 13911 -23 13989 23
rect 14035 -23 14113 23
rect 14159 -23 14237 23
rect 14283 -23 14361 23
rect 14407 -23 14485 23
rect 14531 -23 14609 23
rect 14655 -23 14733 23
rect 14779 -23 14857 23
rect 14903 -23 14981 23
rect 15027 -23 15105 23
rect 15151 -23 15229 23
rect 15275 -23 15353 23
rect 15399 -23 15477 23
rect 15523 -23 15601 23
rect 15647 -23 15725 23
rect 15771 -23 15849 23
rect 15895 -23 15973 23
rect 16019 -23 16097 23
rect 16143 -23 16221 23
rect 16267 -23 16345 23
rect 16391 -23 16469 23
rect 16515 -23 16593 23
rect 16639 -23 16717 23
rect 16763 -23 16841 23
rect 16887 -23 16965 23
rect 17011 -23 17089 23
rect 17135 -23 17213 23
rect 17259 -23 17337 23
rect 17383 -23 17461 23
rect 17507 -23 17585 23
rect 17631 -23 17709 23
rect 17755 -23 17833 23
rect 17879 -23 17957 23
rect 18003 -23 18081 23
rect 18127 -23 18205 23
rect 18251 -23 18329 23
rect 18375 -23 18453 23
rect 18499 -23 18577 23
rect 18623 -23 18701 23
rect 18747 -23 18825 23
rect 18871 -23 18949 23
rect 18995 -23 19073 23
rect 19119 -23 19197 23
rect 19243 -23 19321 23
rect 19367 -23 19445 23
rect 19491 -23 19569 23
rect 19615 -23 19693 23
rect 19739 -23 19817 23
rect 19863 -23 19941 23
rect 19987 -23 20065 23
rect 20111 -23 20189 23
rect 20235 -23 20313 23
rect 20359 -23 20437 23
rect 20483 -23 20561 23
rect 20607 -23 20685 23
rect 20731 -23 20809 23
rect 20855 -23 20933 23
rect 20979 -23 21057 23
rect 21103 -23 21181 23
rect 21227 -23 21305 23
rect 21351 -23 21429 23
rect 21475 -23 21553 23
rect 21599 -23 21677 23
rect 21723 -23 21801 23
rect 21847 -23 21925 23
rect 21971 -23 22049 23
rect 22095 -23 22173 23
rect 22219 -23 22297 23
rect 22343 -23 22421 23
rect 22467 -23 22545 23
rect 22591 -23 22669 23
rect 22715 -23 22793 23
rect 22839 -23 22917 23
rect 22963 -23 23041 23
rect 23087 -23 23165 23
rect 23211 -23 23289 23
rect 23335 -23 23413 23
rect 23459 -23 23537 23
rect 23583 -23 23661 23
rect 23707 -23 23785 23
rect 23831 -23 23909 23
rect 23955 -23 24033 23
rect 24079 -23 24157 23
rect 24203 -23 24281 23
rect 24327 -23 24405 23
rect 24451 -23 24529 23
rect 24575 -23 24653 23
rect 24699 -23 24777 23
rect 24823 -23 24901 23
rect 24947 -23 25025 23
rect 25071 -23 25149 23
rect 25195 -23 25273 23
rect 25319 -23 25397 23
rect 25443 -23 25521 23
rect 25567 -23 25645 23
rect 25691 -23 25769 23
rect 25815 -23 25893 23
rect 25939 -23 26017 23
rect 26063 -23 26141 23
rect 26187 -23 26265 23
rect 26311 -23 26389 23
rect 26435 -23 26513 23
rect 26559 -23 26637 23
rect 26683 -23 26761 23
rect 26807 -23 26885 23
rect 26931 -23 27009 23
rect 27055 -23 27133 23
rect 27179 -23 27257 23
rect 27303 -23 27381 23
rect 27427 -23 27505 23
rect 27551 -23 27629 23
rect 27675 -23 27753 23
rect 27799 -23 27877 23
rect 27923 -23 28001 23
rect 28047 -23 28125 23
rect 28171 -23 28249 23
rect 28295 -23 28373 23
rect 28419 -23 28497 23
rect 28543 -23 28621 23
rect 28667 -23 28745 23
rect 28791 -23 28869 23
rect 28915 -23 28993 23
rect 29039 -23 29117 23
rect 29163 -23 29241 23
rect 29287 -23 29365 23
rect 29411 -23 29489 23
rect 29535 -23 29613 23
rect 29659 -23 29737 23
rect 29783 -23 29861 23
rect 29907 -23 29985 23
rect 30031 -23 30109 23
rect 30155 -23 30233 23
rect 30279 -23 30357 23
rect 30403 -23 30481 23
rect 30527 -23 30605 23
rect 30651 -23 30729 23
rect 30775 -23 30853 23
rect 30899 -23 30977 23
rect 31023 -23 31101 23
rect 31147 -23 31225 23
rect 31271 -23 31349 23
rect 31395 -23 31473 23
rect 31519 -23 31597 23
rect 31643 -23 31721 23
rect 31767 -23 31845 23
rect 31891 -23 31969 23
rect 32015 -23 32093 23
rect 32139 -23 32217 23
rect 32263 -23 32341 23
rect 32387 -23 32465 23
rect 32511 -23 32589 23
rect 32635 -23 32713 23
rect 32759 -23 32837 23
rect 32883 -23 32961 23
rect 33007 -23 33085 23
rect 33131 -23 33209 23
rect 33255 -23 33333 23
rect 33379 -23 33457 23
rect 33503 -23 33581 23
rect 33627 -23 33705 23
rect 33751 -23 33829 23
rect 33875 -23 33953 23
rect 33999 -23 34077 23
rect 34123 -23 34201 23
rect 34247 -23 34325 23
rect 34371 -23 34449 23
rect 34495 -23 34573 23
rect 34619 -23 34697 23
rect 34743 -23 34821 23
rect 34867 -23 34945 23
rect 34991 -23 35069 23
rect 35115 -23 35193 23
rect 35239 -23 35317 23
rect 35363 -23 35441 23
rect 35487 -23 35565 23
rect 35611 -23 35689 23
rect 35735 -23 35813 23
rect 35859 -23 35937 23
rect 35983 -23 36061 23
rect 36107 -23 36185 23
rect 36231 -23 36309 23
rect 36355 -23 36433 23
rect 36479 -23 36557 23
rect 36603 -23 36681 23
rect 36727 -23 36805 23
rect 36851 -23 36929 23
rect 36975 -23 37053 23
rect 37099 -23 37177 23
rect 37223 -23 37301 23
rect 37347 -23 37425 23
rect 37471 -23 37549 23
rect 37595 -23 37673 23
rect 37719 -23 37797 23
rect 37843 -23 37921 23
rect 37967 -23 38045 23
rect 38091 -23 38169 23
rect 38215 -23 38293 23
rect 38339 -23 38417 23
rect 38463 -23 38541 23
rect 38587 -23 38665 23
rect 38711 -23 38789 23
rect 38835 -23 38913 23
rect 38959 -23 39037 23
rect 39083 -23 39161 23
rect 39207 -23 39285 23
rect 39331 -23 39409 23
rect 39455 -23 39533 23
rect 39579 -23 39657 23
rect 39703 -23 39781 23
rect 39827 -23 39905 23
rect 39951 -23 40029 23
rect 40075 -23 40153 23
rect 40199 -23 40277 23
rect 40323 -23 40401 23
rect 40447 -23 40525 23
rect 40571 -23 40649 23
rect 40695 -23 40773 23
rect 40819 -23 40897 23
rect 40943 -23 41021 23
rect 41067 -23 41145 23
rect 41191 -23 41269 23
rect 41315 -23 41393 23
rect 41439 -23 41517 23
rect 41563 -23 41641 23
rect 41687 -23 41765 23
rect 41811 -23 41889 23
rect 41935 -23 42013 23
rect 42059 -23 42137 23
rect 42183 -23 42261 23
rect 42307 -23 42385 23
rect 42431 -23 42509 23
rect 42555 -23 42633 23
rect 42679 -23 42757 23
rect 42803 -23 42881 23
rect 42927 -23 43005 23
rect 43051 -23 43129 23
rect 43175 -23 43253 23
rect 43299 -23 43377 23
rect 43423 -23 43501 23
rect 43547 -23 43625 23
rect 43671 -23 43749 23
rect 43795 -23 43873 23
rect 43919 -23 43997 23
rect 44043 -23 44121 23
rect 44167 -23 44245 23
rect 44291 -23 44369 23
rect 44415 -23 44493 23
rect 44539 -23 44617 23
rect 44663 -23 44741 23
rect 44787 -23 44865 23
rect 44911 -23 44989 23
rect 45035 -23 45113 23
rect 45159 -23 45237 23
rect 45283 -23 45361 23
rect 45407 -23 45485 23
rect 45531 -23 45609 23
rect 45655 -23 45733 23
rect 45779 -23 45857 23
rect 45903 -23 45981 23
rect 46027 -23 46105 23
rect 46151 -23 46229 23
rect 46275 -23 46353 23
rect 46399 -23 46477 23
rect 46523 -23 46601 23
rect 46647 -23 46725 23
rect 46771 -23 46849 23
rect 46895 -23 46973 23
rect 47019 -23 47097 23
rect 47143 -23 47221 23
rect 47267 -23 47345 23
rect 47391 -23 47469 23
rect 47515 -23 47593 23
rect 47639 -23 47717 23
rect 47763 -23 47841 23
rect 47887 -23 47965 23
rect 48011 -23 48089 23
rect 48135 -23 48213 23
rect 48259 -23 48337 23
rect 48383 -23 48461 23
rect 48507 -23 48585 23
rect 48631 -23 48709 23
rect 48755 -23 48833 23
rect 48879 -23 48957 23
rect 49003 -23 49081 23
rect 49127 -23 49205 23
rect 49251 -23 49329 23
rect 49375 -23 49453 23
rect 49499 -23 49577 23
rect 49623 -23 49701 23
rect 49747 -23 49825 23
rect 49871 -23 49949 23
rect 49995 -23 50073 23
rect 50119 -23 50197 23
rect 50243 -23 50321 23
rect 50367 -23 50445 23
rect 50491 -23 50569 23
rect 50615 -23 50693 23
rect 50739 -23 50817 23
rect 50863 -23 50941 23
rect 50987 -23 51065 23
rect 51111 -23 51189 23
rect 51235 -23 51313 23
rect 51359 -23 51437 23
rect 51483 -23 51561 23
rect 51607 -23 51685 23
rect 51731 -23 51809 23
rect 51855 -23 51933 23
rect 51979 -23 52057 23
rect 52103 -23 52181 23
rect 52227 -23 52305 23
rect 52351 -23 52429 23
rect 52475 -23 52553 23
rect 52599 -23 52677 23
rect 52723 -23 52801 23
rect 52847 -23 52925 23
rect 52971 -23 53049 23
rect 53095 -23 53173 23
rect 53219 -23 53297 23
rect 53343 -23 53421 23
rect 53467 -23 53545 23
rect 53591 -23 53669 23
rect 53715 -23 53793 23
rect 53839 -23 53917 23
rect 53963 -23 54041 23
rect 54087 -23 54165 23
rect 54211 -23 54289 23
rect 54335 -23 54413 23
rect 54459 -23 54537 23
rect 54583 -23 54661 23
rect 54707 -23 54785 23
rect 54831 -23 54909 23
rect 54955 -23 55033 23
rect 55079 -23 55157 23
rect 55203 -23 55281 23
rect 55327 -23 55405 23
rect 55451 -23 55529 23
rect 55575 -23 55653 23
rect 55699 -23 55777 23
rect 55823 -23 55901 23
rect 55947 -23 56025 23
rect 56071 -23 56149 23
rect 56195 -23 56273 23
rect 56319 -23 56397 23
rect 56443 -23 56521 23
rect 56567 -23 56645 23
rect 56691 -23 56769 23
rect 56815 -23 56893 23
rect 56939 -23 57017 23
rect 57063 -23 57141 23
rect 57187 -23 57265 23
rect 57311 -23 57389 23
rect 57435 -23 57513 23
rect 57559 -23 57637 23
rect 57683 -23 57761 23
rect 57807 -23 57885 23
rect 57931 -23 58009 23
rect 58055 -23 58133 23
rect 58179 -23 58257 23
rect 58303 -23 58381 23
rect 58427 -23 58505 23
rect 58551 -23 58629 23
rect 58675 -23 58753 23
rect 58799 -23 58877 23
rect 58923 -23 59001 23
rect 59047 -23 59125 23
rect 59171 -23 59249 23
rect 59295 -23 59373 23
rect 59419 -23 59497 23
rect 59543 -23 59621 23
rect 59667 -23 59745 23
rect 59791 -23 59869 23
rect 59915 -23 59993 23
rect 60039 -23 60117 23
rect 60163 -23 60241 23
rect 60287 -23 60365 23
rect 60411 -23 60489 23
rect 60535 -23 60613 23
rect 60659 -23 60737 23
rect 60783 -23 60861 23
rect 60907 -23 60985 23
rect 61031 -23 61109 23
rect 61155 -23 61233 23
rect 61279 -23 61357 23
rect 61403 -23 61481 23
rect 61527 -23 61605 23
rect 61651 -23 61729 23
rect 61775 -23 61853 23
rect 61899 -23 61977 23
rect 62023 -23 62101 23
rect 62147 -23 62225 23
rect 62271 -23 62349 23
rect 62395 -23 62473 23
rect 62519 -23 62597 23
rect 62643 -23 62721 23
rect 62767 -23 62845 23
rect 62891 -23 62969 23
rect 63015 -23 63093 23
rect 63139 -23 63217 23
rect 63263 -23 63341 23
rect 63387 -23 63465 23
rect 63511 -23 63589 23
rect 63635 -23 63713 23
rect 63759 -23 63837 23
rect 63883 -23 63961 23
rect 64007 -23 64085 23
rect 64131 -23 64209 23
rect 64255 -23 64333 23
rect 64379 -23 64457 23
rect 64503 -23 64581 23
rect 64627 -23 64705 23
rect 64751 -23 64829 23
rect 64875 -23 64953 23
rect 64999 -23 65077 23
rect 65123 -23 65201 23
rect 65247 -23 65325 23
rect 65371 -23 65449 23
rect 65495 -23 65573 23
rect 65619 -23 65697 23
rect 65743 -23 65821 23
rect 65867 -23 65945 23
rect 65991 -23 66069 23
rect 66115 -23 66193 23
rect 66239 -23 66317 23
rect 66363 -23 66441 23
rect 66487 -23 66565 23
rect 66611 -23 66689 23
rect 66735 -23 66813 23
rect 66859 -23 66937 23
rect 66983 -23 67061 23
rect 67107 -23 67185 23
rect 67231 -23 67309 23
rect 67355 -23 67433 23
rect 67479 -23 67557 23
rect 67603 -23 67681 23
rect 67727 -23 67805 23
rect 67851 -23 67929 23
rect 67975 -23 68053 23
rect 68099 -23 68177 23
rect 68223 -23 68301 23
rect 68347 -23 68425 23
rect 68471 -23 68549 23
rect 68595 -23 68673 23
rect 68719 -23 68797 23
rect 68843 -23 68921 23
rect 68967 -23 69045 23
rect 69091 -23 69169 23
rect 69215 -23 69293 23
rect 69339 -23 69417 23
rect 69463 -23 69541 23
rect 69587 -23 69665 23
rect 69711 -23 69789 23
rect 69835 -23 69913 23
rect 69959 -23 70037 23
rect 70083 -23 70161 23
rect 70207 -23 70285 23
rect 70331 -23 70409 23
rect 70455 -23 70533 23
rect 70579 -23 70657 23
rect 70703 -23 70781 23
rect 70827 -23 70905 23
rect 70951 -23 71029 23
rect 71075 -23 71153 23
rect 71199 -23 71277 23
rect 71323 -23 71401 23
rect 71447 -23 71525 23
rect 71571 -23 71649 23
rect 71695 -23 71773 23
rect 71819 -23 71897 23
rect 71943 -23 72021 23
rect 72067 -23 72145 23
rect 72191 -23 72269 23
rect 72315 -23 72393 23
rect 72439 -23 72517 23
rect 72563 -23 72641 23
rect 72687 -23 72765 23
rect 72811 -23 72889 23
rect 72935 -23 73013 23
rect 73059 -23 73137 23
rect 73183 -23 73261 23
rect 73307 -23 73385 23
rect 73431 -23 73509 23
rect 73555 -23 73633 23
rect 73679 -23 73757 23
rect 73803 -23 73881 23
rect 73927 -23 74005 23
rect 74051 -23 74129 23
rect 74175 -23 74253 23
rect 74299 -23 74377 23
rect 74423 -23 74501 23
rect 74547 -23 74625 23
rect 74671 -23 74749 23
rect 74795 -23 74873 23
rect 74919 -23 74997 23
rect 75043 -23 75121 23
rect 75167 -23 75245 23
rect 75291 -23 75369 23
rect 75415 -23 75493 23
rect 75539 -23 75617 23
rect 75663 -23 75741 23
rect 75787 -23 75865 23
rect 75911 -23 75989 23
rect 76035 -23 76113 23
rect 76159 -23 76237 23
rect 76283 -23 76361 23
rect 76407 -23 76485 23
rect 76531 -23 76609 23
rect 76655 -23 76733 23
rect 76779 -23 76857 23
rect 76903 -23 76981 23
rect 77027 -23 77105 23
rect 77151 -23 77229 23
rect 77275 -23 77353 23
rect 77399 -23 77477 23
rect 77523 -23 77601 23
rect 77647 -23 77725 23
rect 77771 -23 77849 23
rect 77895 -23 77973 23
rect 78019 -23 78097 23
rect 78143 -23 78221 23
rect 78267 -23 78345 23
rect 78391 -23 78469 23
rect 78515 -23 78593 23
rect 78639 -23 78717 23
rect 78763 -23 78841 23
rect 78887 -23 78965 23
rect 79011 -23 79089 23
rect 79135 -23 79213 23
rect 79259 -23 79337 23
rect 79383 -23 79461 23
rect 79507 -23 79585 23
rect 79631 -23 79709 23
rect 79755 -23 79833 23
rect 79879 -23 79957 23
rect 80003 -23 80081 23
rect 80127 -23 80205 23
rect 80251 -23 80329 23
rect 80375 -23 80453 23
rect 80499 -23 80577 23
rect 80623 -23 80701 23
rect 80747 -23 80825 23
rect 80871 -23 80949 23
rect 80995 -23 81073 23
rect 81119 -23 81197 23
rect 81243 -23 81321 23
rect 81367 -23 81445 23
rect 81491 -23 81569 23
rect 81615 -23 81693 23
rect 81739 -23 81817 23
rect 81863 -23 81941 23
rect 81987 -23 82065 23
rect 82111 -23 82189 23
rect 82235 -23 82313 23
rect 82359 -23 82437 23
rect 82483 -23 82561 23
rect 82607 -23 82685 23
rect 82731 -23 82809 23
rect 82855 -23 82933 23
rect 82979 -23 83057 23
rect 83103 -23 83181 23
rect 83227 -23 83305 23
rect 83351 -23 83429 23
rect 83475 -23 83553 23
rect 83599 -23 83677 23
rect 83723 -23 83801 23
rect 83847 -23 83925 23
rect 83971 -23 84049 23
rect 84095 -23 84173 23
rect 84219 -23 84297 23
rect 84343 -23 84421 23
rect 84467 -23 84545 23
rect 84591 -23 84669 23
rect 84715 -23 84793 23
rect 84839 -23 84917 23
rect 84963 -23 85041 23
rect 85087 -23 85165 23
rect 85211 -23 85289 23
rect 85335 -23 85413 23
rect 85459 -23 85537 23
rect 85583 -23 85602 23
rect -42 -42 85602 -23
<< psubdiffcont >>
rect -23 349 23 395
rect 101 349 147 395
rect 225 349 271 395
rect 349 349 395 395
rect 473 349 519 395
rect 597 349 643 395
rect 721 349 767 395
rect 845 349 891 395
rect 969 349 1015 395
rect 1093 349 1139 395
rect 1217 349 1263 395
rect 1341 349 1387 395
rect 1465 349 1511 395
rect 1589 349 1635 395
rect 1713 349 1759 395
rect 1837 349 1883 395
rect 1961 349 2007 395
rect 2085 349 2131 395
rect 2209 349 2255 395
rect 2333 349 2379 395
rect 2457 349 2503 395
rect 2581 349 2627 395
rect 2705 349 2751 395
rect 2829 349 2875 395
rect 2953 349 2999 395
rect 3077 349 3123 395
rect 3201 349 3247 395
rect 3325 349 3371 395
rect 3449 349 3495 395
rect 3573 349 3619 395
rect 3697 349 3743 395
rect 3821 349 3867 395
rect 3945 349 3991 395
rect 4069 349 4115 395
rect 4193 349 4239 395
rect 4317 349 4363 395
rect 4441 349 4487 395
rect 4565 349 4611 395
rect 4689 349 4735 395
rect 4813 349 4859 395
rect 4937 349 4983 395
rect 5061 349 5107 395
rect 5185 349 5231 395
rect 5309 349 5355 395
rect 5433 349 5479 395
rect 5557 349 5603 395
rect 5681 349 5727 395
rect 5805 349 5851 395
rect 5929 349 5975 395
rect 6053 349 6099 395
rect 6177 349 6223 395
rect 6301 349 6347 395
rect 6425 349 6471 395
rect 6549 349 6595 395
rect 6673 349 6719 395
rect 6797 349 6843 395
rect 6921 349 6967 395
rect 7045 349 7091 395
rect 7169 349 7215 395
rect 7293 349 7339 395
rect 7417 349 7463 395
rect 7541 349 7587 395
rect 7665 349 7711 395
rect 7789 349 7835 395
rect 7913 349 7959 395
rect 8037 349 8083 395
rect 8161 349 8207 395
rect 8285 349 8331 395
rect 8409 349 8455 395
rect 8533 349 8579 395
rect 8657 349 8703 395
rect 8781 349 8827 395
rect 8905 349 8951 395
rect 9029 349 9075 395
rect 9153 349 9199 395
rect 9277 349 9323 395
rect 9401 349 9447 395
rect 9525 349 9571 395
rect 9649 349 9695 395
rect 9773 349 9819 395
rect 9897 349 9943 395
rect 10021 349 10067 395
rect 10145 349 10191 395
rect 10269 349 10315 395
rect 10393 349 10439 395
rect 10517 349 10563 395
rect 10641 349 10687 395
rect 10765 349 10811 395
rect 10889 349 10935 395
rect 11013 349 11059 395
rect 11137 349 11183 395
rect 11261 349 11307 395
rect 11385 349 11431 395
rect 11509 349 11555 395
rect 11633 349 11679 395
rect 11757 349 11803 395
rect 11881 349 11927 395
rect 12005 349 12051 395
rect 12129 349 12175 395
rect 12253 349 12299 395
rect 12377 349 12423 395
rect 12501 349 12547 395
rect 12625 349 12671 395
rect 12749 349 12795 395
rect 12873 349 12919 395
rect 12997 349 13043 395
rect 13121 349 13167 395
rect 13245 349 13291 395
rect 13369 349 13415 395
rect 13493 349 13539 395
rect 13617 349 13663 395
rect 13741 349 13787 395
rect 13865 349 13911 395
rect 13989 349 14035 395
rect 14113 349 14159 395
rect 14237 349 14283 395
rect 14361 349 14407 395
rect 14485 349 14531 395
rect 14609 349 14655 395
rect 14733 349 14779 395
rect 14857 349 14903 395
rect 14981 349 15027 395
rect 15105 349 15151 395
rect 15229 349 15275 395
rect 15353 349 15399 395
rect 15477 349 15523 395
rect 15601 349 15647 395
rect 15725 349 15771 395
rect 15849 349 15895 395
rect 15973 349 16019 395
rect 16097 349 16143 395
rect 16221 349 16267 395
rect 16345 349 16391 395
rect 16469 349 16515 395
rect 16593 349 16639 395
rect 16717 349 16763 395
rect 16841 349 16887 395
rect 16965 349 17011 395
rect 17089 349 17135 395
rect 17213 349 17259 395
rect 17337 349 17383 395
rect 17461 349 17507 395
rect 17585 349 17631 395
rect 17709 349 17755 395
rect 17833 349 17879 395
rect 17957 349 18003 395
rect 18081 349 18127 395
rect 18205 349 18251 395
rect 18329 349 18375 395
rect 18453 349 18499 395
rect 18577 349 18623 395
rect 18701 349 18747 395
rect 18825 349 18871 395
rect 18949 349 18995 395
rect 19073 349 19119 395
rect 19197 349 19243 395
rect 19321 349 19367 395
rect 19445 349 19491 395
rect 19569 349 19615 395
rect 19693 349 19739 395
rect 19817 349 19863 395
rect 19941 349 19987 395
rect 20065 349 20111 395
rect 20189 349 20235 395
rect 20313 349 20359 395
rect 20437 349 20483 395
rect 20561 349 20607 395
rect 20685 349 20731 395
rect 20809 349 20855 395
rect 20933 349 20979 395
rect 21057 349 21103 395
rect 21181 349 21227 395
rect 21305 349 21351 395
rect 21429 349 21475 395
rect 21553 349 21599 395
rect 21677 349 21723 395
rect 21801 349 21847 395
rect 21925 349 21971 395
rect 22049 349 22095 395
rect 22173 349 22219 395
rect 22297 349 22343 395
rect 22421 349 22467 395
rect 22545 349 22591 395
rect 22669 349 22715 395
rect 22793 349 22839 395
rect 22917 349 22963 395
rect 23041 349 23087 395
rect 23165 349 23211 395
rect 23289 349 23335 395
rect 23413 349 23459 395
rect 23537 349 23583 395
rect 23661 349 23707 395
rect 23785 349 23831 395
rect 23909 349 23955 395
rect 24033 349 24079 395
rect 24157 349 24203 395
rect 24281 349 24327 395
rect 24405 349 24451 395
rect 24529 349 24575 395
rect 24653 349 24699 395
rect 24777 349 24823 395
rect 24901 349 24947 395
rect 25025 349 25071 395
rect 25149 349 25195 395
rect 25273 349 25319 395
rect 25397 349 25443 395
rect 25521 349 25567 395
rect 25645 349 25691 395
rect 25769 349 25815 395
rect 25893 349 25939 395
rect 26017 349 26063 395
rect 26141 349 26187 395
rect 26265 349 26311 395
rect 26389 349 26435 395
rect 26513 349 26559 395
rect 26637 349 26683 395
rect 26761 349 26807 395
rect 26885 349 26931 395
rect 27009 349 27055 395
rect 27133 349 27179 395
rect 27257 349 27303 395
rect 27381 349 27427 395
rect 27505 349 27551 395
rect 27629 349 27675 395
rect 27753 349 27799 395
rect 27877 349 27923 395
rect 28001 349 28047 395
rect 28125 349 28171 395
rect 28249 349 28295 395
rect 28373 349 28419 395
rect 28497 349 28543 395
rect 28621 349 28667 395
rect 28745 349 28791 395
rect 28869 349 28915 395
rect 28993 349 29039 395
rect 29117 349 29163 395
rect 29241 349 29287 395
rect 29365 349 29411 395
rect 29489 349 29535 395
rect 29613 349 29659 395
rect 29737 349 29783 395
rect 29861 349 29907 395
rect 29985 349 30031 395
rect 30109 349 30155 395
rect 30233 349 30279 395
rect 30357 349 30403 395
rect 30481 349 30527 395
rect 30605 349 30651 395
rect 30729 349 30775 395
rect 30853 349 30899 395
rect 30977 349 31023 395
rect 31101 349 31147 395
rect 31225 349 31271 395
rect 31349 349 31395 395
rect 31473 349 31519 395
rect 31597 349 31643 395
rect 31721 349 31767 395
rect 31845 349 31891 395
rect 31969 349 32015 395
rect 32093 349 32139 395
rect 32217 349 32263 395
rect 32341 349 32387 395
rect 32465 349 32511 395
rect 32589 349 32635 395
rect 32713 349 32759 395
rect 32837 349 32883 395
rect 32961 349 33007 395
rect 33085 349 33131 395
rect 33209 349 33255 395
rect 33333 349 33379 395
rect 33457 349 33503 395
rect 33581 349 33627 395
rect 33705 349 33751 395
rect 33829 349 33875 395
rect 33953 349 33999 395
rect 34077 349 34123 395
rect 34201 349 34247 395
rect 34325 349 34371 395
rect 34449 349 34495 395
rect 34573 349 34619 395
rect 34697 349 34743 395
rect 34821 349 34867 395
rect 34945 349 34991 395
rect 35069 349 35115 395
rect 35193 349 35239 395
rect 35317 349 35363 395
rect 35441 349 35487 395
rect 35565 349 35611 395
rect 35689 349 35735 395
rect 35813 349 35859 395
rect 35937 349 35983 395
rect 36061 349 36107 395
rect 36185 349 36231 395
rect 36309 349 36355 395
rect 36433 349 36479 395
rect 36557 349 36603 395
rect 36681 349 36727 395
rect 36805 349 36851 395
rect 36929 349 36975 395
rect 37053 349 37099 395
rect 37177 349 37223 395
rect 37301 349 37347 395
rect 37425 349 37471 395
rect 37549 349 37595 395
rect 37673 349 37719 395
rect 37797 349 37843 395
rect 37921 349 37967 395
rect 38045 349 38091 395
rect 38169 349 38215 395
rect 38293 349 38339 395
rect 38417 349 38463 395
rect 38541 349 38587 395
rect 38665 349 38711 395
rect 38789 349 38835 395
rect 38913 349 38959 395
rect 39037 349 39083 395
rect 39161 349 39207 395
rect 39285 349 39331 395
rect 39409 349 39455 395
rect 39533 349 39579 395
rect 39657 349 39703 395
rect 39781 349 39827 395
rect 39905 349 39951 395
rect 40029 349 40075 395
rect 40153 349 40199 395
rect 40277 349 40323 395
rect 40401 349 40447 395
rect 40525 349 40571 395
rect 40649 349 40695 395
rect 40773 349 40819 395
rect 40897 349 40943 395
rect 41021 349 41067 395
rect 41145 349 41191 395
rect 41269 349 41315 395
rect 41393 349 41439 395
rect 41517 349 41563 395
rect 41641 349 41687 395
rect 41765 349 41811 395
rect 41889 349 41935 395
rect 42013 349 42059 395
rect 42137 349 42183 395
rect 42261 349 42307 395
rect 42385 349 42431 395
rect 42509 349 42555 395
rect 42633 349 42679 395
rect 42757 349 42803 395
rect 42881 349 42927 395
rect 43005 349 43051 395
rect 43129 349 43175 395
rect 43253 349 43299 395
rect 43377 349 43423 395
rect 43501 349 43547 395
rect 43625 349 43671 395
rect 43749 349 43795 395
rect 43873 349 43919 395
rect 43997 349 44043 395
rect 44121 349 44167 395
rect 44245 349 44291 395
rect 44369 349 44415 395
rect 44493 349 44539 395
rect 44617 349 44663 395
rect 44741 349 44787 395
rect 44865 349 44911 395
rect 44989 349 45035 395
rect 45113 349 45159 395
rect 45237 349 45283 395
rect 45361 349 45407 395
rect 45485 349 45531 395
rect 45609 349 45655 395
rect 45733 349 45779 395
rect 45857 349 45903 395
rect 45981 349 46027 395
rect 46105 349 46151 395
rect 46229 349 46275 395
rect 46353 349 46399 395
rect 46477 349 46523 395
rect 46601 349 46647 395
rect 46725 349 46771 395
rect 46849 349 46895 395
rect 46973 349 47019 395
rect 47097 349 47143 395
rect 47221 349 47267 395
rect 47345 349 47391 395
rect 47469 349 47515 395
rect 47593 349 47639 395
rect 47717 349 47763 395
rect 47841 349 47887 395
rect 47965 349 48011 395
rect 48089 349 48135 395
rect 48213 349 48259 395
rect 48337 349 48383 395
rect 48461 349 48507 395
rect 48585 349 48631 395
rect 48709 349 48755 395
rect 48833 349 48879 395
rect 48957 349 49003 395
rect 49081 349 49127 395
rect 49205 349 49251 395
rect 49329 349 49375 395
rect 49453 349 49499 395
rect 49577 349 49623 395
rect 49701 349 49747 395
rect 49825 349 49871 395
rect 49949 349 49995 395
rect 50073 349 50119 395
rect 50197 349 50243 395
rect 50321 349 50367 395
rect 50445 349 50491 395
rect 50569 349 50615 395
rect 50693 349 50739 395
rect 50817 349 50863 395
rect 50941 349 50987 395
rect 51065 349 51111 395
rect 51189 349 51235 395
rect 51313 349 51359 395
rect 51437 349 51483 395
rect 51561 349 51607 395
rect 51685 349 51731 395
rect 51809 349 51855 395
rect 51933 349 51979 395
rect 52057 349 52103 395
rect 52181 349 52227 395
rect 52305 349 52351 395
rect 52429 349 52475 395
rect 52553 349 52599 395
rect 52677 349 52723 395
rect 52801 349 52847 395
rect 52925 349 52971 395
rect 53049 349 53095 395
rect 53173 349 53219 395
rect 53297 349 53343 395
rect 53421 349 53467 395
rect 53545 349 53591 395
rect 53669 349 53715 395
rect 53793 349 53839 395
rect 53917 349 53963 395
rect 54041 349 54087 395
rect 54165 349 54211 395
rect 54289 349 54335 395
rect 54413 349 54459 395
rect 54537 349 54583 395
rect 54661 349 54707 395
rect 54785 349 54831 395
rect 54909 349 54955 395
rect 55033 349 55079 395
rect 55157 349 55203 395
rect 55281 349 55327 395
rect 55405 349 55451 395
rect 55529 349 55575 395
rect 55653 349 55699 395
rect 55777 349 55823 395
rect 55901 349 55947 395
rect 56025 349 56071 395
rect 56149 349 56195 395
rect 56273 349 56319 395
rect 56397 349 56443 395
rect 56521 349 56567 395
rect 56645 349 56691 395
rect 56769 349 56815 395
rect 56893 349 56939 395
rect 57017 349 57063 395
rect 57141 349 57187 395
rect 57265 349 57311 395
rect 57389 349 57435 395
rect 57513 349 57559 395
rect 57637 349 57683 395
rect 57761 349 57807 395
rect 57885 349 57931 395
rect 58009 349 58055 395
rect 58133 349 58179 395
rect 58257 349 58303 395
rect 58381 349 58427 395
rect 58505 349 58551 395
rect 58629 349 58675 395
rect 58753 349 58799 395
rect 58877 349 58923 395
rect 59001 349 59047 395
rect 59125 349 59171 395
rect 59249 349 59295 395
rect 59373 349 59419 395
rect 59497 349 59543 395
rect 59621 349 59667 395
rect 59745 349 59791 395
rect 59869 349 59915 395
rect 59993 349 60039 395
rect 60117 349 60163 395
rect 60241 349 60287 395
rect 60365 349 60411 395
rect 60489 349 60535 395
rect 60613 349 60659 395
rect 60737 349 60783 395
rect 60861 349 60907 395
rect 60985 349 61031 395
rect 61109 349 61155 395
rect 61233 349 61279 395
rect 61357 349 61403 395
rect 61481 349 61527 395
rect 61605 349 61651 395
rect 61729 349 61775 395
rect 61853 349 61899 395
rect 61977 349 62023 395
rect 62101 349 62147 395
rect 62225 349 62271 395
rect 62349 349 62395 395
rect 62473 349 62519 395
rect 62597 349 62643 395
rect 62721 349 62767 395
rect 62845 349 62891 395
rect 62969 349 63015 395
rect 63093 349 63139 395
rect 63217 349 63263 395
rect 63341 349 63387 395
rect 63465 349 63511 395
rect 63589 349 63635 395
rect 63713 349 63759 395
rect 63837 349 63883 395
rect 63961 349 64007 395
rect 64085 349 64131 395
rect 64209 349 64255 395
rect 64333 349 64379 395
rect 64457 349 64503 395
rect 64581 349 64627 395
rect 64705 349 64751 395
rect 64829 349 64875 395
rect 64953 349 64999 395
rect 65077 349 65123 395
rect 65201 349 65247 395
rect 65325 349 65371 395
rect 65449 349 65495 395
rect 65573 349 65619 395
rect 65697 349 65743 395
rect 65821 349 65867 395
rect 65945 349 65991 395
rect 66069 349 66115 395
rect 66193 349 66239 395
rect 66317 349 66363 395
rect 66441 349 66487 395
rect 66565 349 66611 395
rect 66689 349 66735 395
rect 66813 349 66859 395
rect 66937 349 66983 395
rect 67061 349 67107 395
rect 67185 349 67231 395
rect 67309 349 67355 395
rect 67433 349 67479 395
rect 67557 349 67603 395
rect 67681 349 67727 395
rect 67805 349 67851 395
rect 67929 349 67975 395
rect 68053 349 68099 395
rect 68177 349 68223 395
rect 68301 349 68347 395
rect 68425 349 68471 395
rect 68549 349 68595 395
rect 68673 349 68719 395
rect 68797 349 68843 395
rect 68921 349 68967 395
rect 69045 349 69091 395
rect 69169 349 69215 395
rect 69293 349 69339 395
rect 69417 349 69463 395
rect 69541 349 69587 395
rect 69665 349 69711 395
rect 69789 349 69835 395
rect 69913 349 69959 395
rect 70037 349 70083 395
rect 70161 349 70207 395
rect 70285 349 70331 395
rect 70409 349 70455 395
rect 70533 349 70579 395
rect 70657 349 70703 395
rect 70781 349 70827 395
rect 70905 349 70951 395
rect 71029 349 71075 395
rect 71153 349 71199 395
rect 71277 349 71323 395
rect 71401 349 71447 395
rect 71525 349 71571 395
rect 71649 349 71695 395
rect 71773 349 71819 395
rect 71897 349 71943 395
rect 72021 349 72067 395
rect 72145 349 72191 395
rect 72269 349 72315 395
rect 72393 349 72439 395
rect 72517 349 72563 395
rect 72641 349 72687 395
rect 72765 349 72811 395
rect 72889 349 72935 395
rect 73013 349 73059 395
rect 73137 349 73183 395
rect 73261 349 73307 395
rect 73385 349 73431 395
rect 73509 349 73555 395
rect 73633 349 73679 395
rect 73757 349 73803 395
rect 73881 349 73927 395
rect 74005 349 74051 395
rect 74129 349 74175 395
rect 74253 349 74299 395
rect 74377 349 74423 395
rect 74501 349 74547 395
rect 74625 349 74671 395
rect 74749 349 74795 395
rect 74873 349 74919 395
rect 74997 349 75043 395
rect 75121 349 75167 395
rect 75245 349 75291 395
rect 75369 349 75415 395
rect 75493 349 75539 395
rect 75617 349 75663 395
rect 75741 349 75787 395
rect 75865 349 75911 395
rect 75989 349 76035 395
rect 76113 349 76159 395
rect 76237 349 76283 395
rect 76361 349 76407 395
rect 76485 349 76531 395
rect 76609 349 76655 395
rect 76733 349 76779 395
rect 76857 349 76903 395
rect 76981 349 77027 395
rect 77105 349 77151 395
rect 77229 349 77275 395
rect 77353 349 77399 395
rect 77477 349 77523 395
rect 77601 349 77647 395
rect 77725 349 77771 395
rect 77849 349 77895 395
rect 77973 349 78019 395
rect 78097 349 78143 395
rect 78221 349 78267 395
rect 78345 349 78391 395
rect 78469 349 78515 395
rect 78593 349 78639 395
rect 78717 349 78763 395
rect 78841 349 78887 395
rect 78965 349 79011 395
rect 79089 349 79135 395
rect 79213 349 79259 395
rect 79337 349 79383 395
rect 79461 349 79507 395
rect 79585 349 79631 395
rect 79709 349 79755 395
rect 79833 349 79879 395
rect 79957 349 80003 395
rect 80081 349 80127 395
rect 80205 349 80251 395
rect 80329 349 80375 395
rect 80453 349 80499 395
rect 80577 349 80623 395
rect 80701 349 80747 395
rect 80825 349 80871 395
rect 80949 349 80995 395
rect 81073 349 81119 395
rect 81197 349 81243 395
rect 81321 349 81367 395
rect 81445 349 81491 395
rect 81569 349 81615 395
rect 81693 349 81739 395
rect 81817 349 81863 395
rect 81941 349 81987 395
rect 82065 349 82111 395
rect 82189 349 82235 395
rect 82313 349 82359 395
rect 82437 349 82483 395
rect 82561 349 82607 395
rect 82685 349 82731 395
rect 82809 349 82855 395
rect 82933 349 82979 395
rect 83057 349 83103 395
rect 83181 349 83227 395
rect 83305 349 83351 395
rect 83429 349 83475 395
rect 83553 349 83599 395
rect 83677 349 83723 395
rect 83801 349 83847 395
rect 83925 349 83971 395
rect 84049 349 84095 395
rect 84173 349 84219 395
rect 84297 349 84343 395
rect 84421 349 84467 395
rect 84545 349 84591 395
rect 84669 349 84715 395
rect 84793 349 84839 395
rect 84917 349 84963 395
rect 85041 349 85087 395
rect 85165 349 85211 395
rect 85289 349 85335 395
rect 85413 349 85459 395
rect 85537 349 85583 395
rect -23 225 23 271
rect 101 225 147 271
rect 225 225 271 271
rect 349 225 395 271
rect 473 225 519 271
rect 597 225 643 271
rect 721 225 767 271
rect 845 225 891 271
rect 969 225 1015 271
rect 1093 225 1139 271
rect 1217 225 1263 271
rect 1341 225 1387 271
rect 1465 225 1511 271
rect 1589 225 1635 271
rect 1713 225 1759 271
rect 1837 225 1883 271
rect 1961 225 2007 271
rect 2085 225 2131 271
rect 2209 225 2255 271
rect 2333 225 2379 271
rect 2457 225 2503 271
rect 2581 225 2627 271
rect 2705 225 2751 271
rect 2829 225 2875 271
rect 2953 225 2999 271
rect 3077 225 3123 271
rect 3201 225 3247 271
rect 3325 225 3371 271
rect 3449 225 3495 271
rect 3573 225 3619 271
rect 3697 225 3743 271
rect 3821 225 3867 271
rect 3945 225 3991 271
rect 4069 225 4115 271
rect 4193 225 4239 271
rect 4317 225 4363 271
rect 4441 225 4487 271
rect 4565 225 4611 271
rect 4689 225 4735 271
rect 4813 225 4859 271
rect 4937 225 4983 271
rect 5061 225 5107 271
rect 5185 225 5231 271
rect 5309 225 5355 271
rect 5433 225 5479 271
rect 5557 225 5603 271
rect 5681 225 5727 271
rect 5805 225 5851 271
rect 5929 225 5975 271
rect 6053 225 6099 271
rect 6177 225 6223 271
rect 6301 225 6347 271
rect 6425 225 6471 271
rect 6549 225 6595 271
rect 6673 225 6719 271
rect 6797 225 6843 271
rect 6921 225 6967 271
rect 7045 225 7091 271
rect 7169 225 7215 271
rect 7293 225 7339 271
rect 7417 225 7463 271
rect 7541 225 7587 271
rect 7665 225 7711 271
rect 7789 225 7835 271
rect 7913 225 7959 271
rect 8037 225 8083 271
rect 8161 225 8207 271
rect 8285 225 8331 271
rect 8409 225 8455 271
rect 8533 225 8579 271
rect 8657 225 8703 271
rect 8781 225 8827 271
rect 8905 225 8951 271
rect 9029 225 9075 271
rect 9153 225 9199 271
rect 9277 225 9323 271
rect 9401 225 9447 271
rect 9525 225 9571 271
rect 9649 225 9695 271
rect 9773 225 9819 271
rect 9897 225 9943 271
rect 10021 225 10067 271
rect 10145 225 10191 271
rect 10269 225 10315 271
rect 10393 225 10439 271
rect 10517 225 10563 271
rect 10641 225 10687 271
rect 10765 225 10811 271
rect 10889 225 10935 271
rect 11013 225 11059 271
rect 11137 225 11183 271
rect 11261 225 11307 271
rect 11385 225 11431 271
rect 11509 225 11555 271
rect 11633 225 11679 271
rect 11757 225 11803 271
rect 11881 225 11927 271
rect 12005 225 12051 271
rect 12129 225 12175 271
rect 12253 225 12299 271
rect 12377 225 12423 271
rect 12501 225 12547 271
rect 12625 225 12671 271
rect 12749 225 12795 271
rect 12873 225 12919 271
rect 12997 225 13043 271
rect 13121 225 13167 271
rect 13245 225 13291 271
rect 13369 225 13415 271
rect 13493 225 13539 271
rect 13617 225 13663 271
rect 13741 225 13787 271
rect 13865 225 13911 271
rect 13989 225 14035 271
rect 14113 225 14159 271
rect 14237 225 14283 271
rect 14361 225 14407 271
rect 14485 225 14531 271
rect 14609 225 14655 271
rect 14733 225 14779 271
rect 14857 225 14903 271
rect 14981 225 15027 271
rect 15105 225 15151 271
rect 15229 225 15275 271
rect 15353 225 15399 271
rect 15477 225 15523 271
rect 15601 225 15647 271
rect 15725 225 15771 271
rect 15849 225 15895 271
rect 15973 225 16019 271
rect 16097 225 16143 271
rect 16221 225 16267 271
rect 16345 225 16391 271
rect 16469 225 16515 271
rect 16593 225 16639 271
rect 16717 225 16763 271
rect 16841 225 16887 271
rect 16965 225 17011 271
rect 17089 225 17135 271
rect 17213 225 17259 271
rect 17337 225 17383 271
rect 17461 225 17507 271
rect 17585 225 17631 271
rect 17709 225 17755 271
rect 17833 225 17879 271
rect 17957 225 18003 271
rect 18081 225 18127 271
rect 18205 225 18251 271
rect 18329 225 18375 271
rect 18453 225 18499 271
rect 18577 225 18623 271
rect 18701 225 18747 271
rect 18825 225 18871 271
rect 18949 225 18995 271
rect 19073 225 19119 271
rect 19197 225 19243 271
rect 19321 225 19367 271
rect 19445 225 19491 271
rect 19569 225 19615 271
rect 19693 225 19739 271
rect 19817 225 19863 271
rect 19941 225 19987 271
rect 20065 225 20111 271
rect 20189 225 20235 271
rect 20313 225 20359 271
rect 20437 225 20483 271
rect 20561 225 20607 271
rect 20685 225 20731 271
rect 20809 225 20855 271
rect 20933 225 20979 271
rect 21057 225 21103 271
rect 21181 225 21227 271
rect 21305 225 21351 271
rect 21429 225 21475 271
rect 21553 225 21599 271
rect 21677 225 21723 271
rect 21801 225 21847 271
rect 21925 225 21971 271
rect 22049 225 22095 271
rect 22173 225 22219 271
rect 22297 225 22343 271
rect 22421 225 22467 271
rect 22545 225 22591 271
rect 22669 225 22715 271
rect 22793 225 22839 271
rect 22917 225 22963 271
rect 23041 225 23087 271
rect 23165 225 23211 271
rect 23289 225 23335 271
rect 23413 225 23459 271
rect 23537 225 23583 271
rect 23661 225 23707 271
rect 23785 225 23831 271
rect 23909 225 23955 271
rect 24033 225 24079 271
rect 24157 225 24203 271
rect 24281 225 24327 271
rect 24405 225 24451 271
rect 24529 225 24575 271
rect 24653 225 24699 271
rect 24777 225 24823 271
rect 24901 225 24947 271
rect 25025 225 25071 271
rect 25149 225 25195 271
rect 25273 225 25319 271
rect 25397 225 25443 271
rect 25521 225 25567 271
rect 25645 225 25691 271
rect 25769 225 25815 271
rect 25893 225 25939 271
rect 26017 225 26063 271
rect 26141 225 26187 271
rect 26265 225 26311 271
rect 26389 225 26435 271
rect 26513 225 26559 271
rect 26637 225 26683 271
rect 26761 225 26807 271
rect 26885 225 26931 271
rect 27009 225 27055 271
rect 27133 225 27179 271
rect 27257 225 27303 271
rect 27381 225 27427 271
rect 27505 225 27551 271
rect 27629 225 27675 271
rect 27753 225 27799 271
rect 27877 225 27923 271
rect 28001 225 28047 271
rect 28125 225 28171 271
rect 28249 225 28295 271
rect 28373 225 28419 271
rect 28497 225 28543 271
rect 28621 225 28667 271
rect 28745 225 28791 271
rect 28869 225 28915 271
rect 28993 225 29039 271
rect 29117 225 29163 271
rect 29241 225 29287 271
rect 29365 225 29411 271
rect 29489 225 29535 271
rect 29613 225 29659 271
rect 29737 225 29783 271
rect 29861 225 29907 271
rect 29985 225 30031 271
rect 30109 225 30155 271
rect 30233 225 30279 271
rect 30357 225 30403 271
rect 30481 225 30527 271
rect 30605 225 30651 271
rect 30729 225 30775 271
rect 30853 225 30899 271
rect 30977 225 31023 271
rect 31101 225 31147 271
rect 31225 225 31271 271
rect 31349 225 31395 271
rect 31473 225 31519 271
rect 31597 225 31643 271
rect 31721 225 31767 271
rect 31845 225 31891 271
rect 31969 225 32015 271
rect 32093 225 32139 271
rect 32217 225 32263 271
rect 32341 225 32387 271
rect 32465 225 32511 271
rect 32589 225 32635 271
rect 32713 225 32759 271
rect 32837 225 32883 271
rect 32961 225 33007 271
rect 33085 225 33131 271
rect 33209 225 33255 271
rect 33333 225 33379 271
rect 33457 225 33503 271
rect 33581 225 33627 271
rect 33705 225 33751 271
rect 33829 225 33875 271
rect 33953 225 33999 271
rect 34077 225 34123 271
rect 34201 225 34247 271
rect 34325 225 34371 271
rect 34449 225 34495 271
rect 34573 225 34619 271
rect 34697 225 34743 271
rect 34821 225 34867 271
rect 34945 225 34991 271
rect 35069 225 35115 271
rect 35193 225 35239 271
rect 35317 225 35363 271
rect 35441 225 35487 271
rect 35565 225 35611 271
rect 35689 225 35735 271
rect 35813 225 35859 271
rect 35937 225 35983 271
rect 36061 225 36107 271
rect 36185 225 36231 271
rect 36309 225 36355 271
rect 36433 225 36479 271
rect 36557 225 36603 271
rect 36681 225 36727 271
rect 36805 225 36851 271
rect 36929 225 36975 271
rect 37053 225 37099 271
rect 37177 225 37223 271
rect 37301 225 37347 271
rect 37425 225 37471 271
rect 37549 225 37595 271
rect 37673 225 37719 271
rect 37797 225 37843 271
rect 37921 225 37967 271
rect 38045 225 38091 271
rect 38169 225 38215 271
rect 38293 225 38339 271
rect 38417 225 38463 271
rect 38541 225 38587 271
rect 38665 225 38711 271
rect 38789 225 38835 271
rect 38913 225 38959 271
rect 39037 225 39083 271
rect 39161 225 39207 271
rect 39285 225 39331 271
rect 39409 225 39455 271
rect 39533 225 39579 271
rect 39657 225 39703 271
rect 39781 225 39827 271
rect 39905 225 39951 271
rect 40029 225 40075 271
rect 40153 225 40199 271
rect 40277 225 40323 271
rect 40401 225 40447 271
rect 40525 225 40571 271
rect 40649 225 40695 271
rect 40773 225 40819 271
rect 40897 225 40943 271
rect 41021 225 41067 271
rect 41145 225 41191 271
rect 41269 225 41315 271
rect 41393 225 41439 271
rect 41517 225 41563 271
rect 41641 225 41687 271
rect 41765 225 41811 271
rect 41889 225 41935 271
rect 42013 225 42059 271
rect 42137 225 42183 271
rect 42261 225 42307 271
rect 42385 225 42431 271
rect 42509 225 42555 271
rect 42633 225 42679 271
rect 42757 225 42803 271
rect 42881 225 42927 271
rect 43005 225 43051 271
rect 43129 225 43175 271
rect 43253 225 43299 271
rect 43377 225 43423 271
rect 43501 225 43547 271
rect 43625 225 43671 271
rect 43749 225 43795 271
rect 43873 225 43919 271
rect 43997 225 44043 271
rect 44121 225 44167 271
rect 44245 225 44291 271
rect 44369 225 44415 271
rect 44493 225 44539 271
rect 44617 225 44663 271
rect 44741 225 44787 271
rect 44865 225 44911 271
rect 44989 225 45035 271
rect 45113 225 45159 271
rect 45237 225 45283 271
rect 45361 225 45407 271
rect 45485 225 45531 271
rect 45609 225 45655 271
rect 45733 225 45779 271
rect 45857 225 45903 271
rect 45981 225 46027 271
rect 46105 225 46151 271
rect 46229 225 46275 271
rect 46353 225 46399 271
rect 46477 225 46523 271
rect 46601 225 46647 271
rect 46725 225 46771 271
rect 46849 225 46895 271
rect 46973 225 47019 271
rect 47097 225 47143 271
rect 47221 225 47267 271
rect 47345 225 47391 271
rect 47469 225 47515 271
rect 47593 225 47639 271
rect 47717 225 47763 271
rect 47841 225 47887 271
rect 47965 225 48011 271
rect 48089 225 48135 271
rect 48213 225 48259 271
rect 48337 225 48383 271
rect 48461 225 48507 271
rect 48585 225 48631 271
rect 48709 225 48755 271
rect 48833 225 48879 271
rect 48957 225 49003 271
rect 49081 225 49127 271
rect 49205 225 49251 271
rect 49329 225 49375 271
rect 49453 225 49499 271
rect 49577 225 49623 271
rect 49701 225 49747 271
rect 49825 225 49871 271
rect 49949 225 49995 271
rect 50073 225 50119 271
rect 50197 225 50243 271
rect 50321 225 50367 271
rect 50445 225 50491 271
rect 50569 225 50615 271
rect 50693 225 50739 271
rect 50817 225 50863 271
rect 50941 225 50987 271
rect 51065 225 51111 271
rect 51189 225 51235 271
rect 51313 225 51359 271
rect 51437 225 51483 271
rect 51561 225 51607 271
rect 51685 225 51731 271
rect 51809 225 51855 271
rect 51933 225 51979 271
rect 52057 225 52103 271
rect 52181 225 52227 271
rect 52305 225 52351 271
rect 52429 225 52475 271
rect 52553 225 52599 271
rect 52677 225 52723 271
rect 52801 225 52847 271
rect 52925 225 52971 271
rect 53049 225 53095 271
rect 53173 225 53219 271
rect 53297 225 53343 271
rect 53421 225 53467 271
rect 53545 225 53591 271
rect 53669 225 53715 271
rect 53793 225 53839 271
rect 53917 225 53963 271
rect 54041 225 54087 271
rect 54165 225 54211 271
rect 54289 225 54335 271
rect 54413 225 54459 271
rect 54537 225 54583 271
rect 54661 225 54707 271
rect 54785 225 54831 271
rect 54909 225 54955 271
rect 55033 225 55079 271
rect 55157 225 55203 271
rect 55281 225 55327 271
rect 55405 225 55451 271
rect 55529 225 55575 271
rect 55653 225 55699 271
rect 55777 225 55823 271
rect 55901 225 55947 271
rect 56025 225 56071 271
rect 56149 225 56195 271
rect 56273 225 56319 271
rect 56397 225 56443 271
rect 56521 225 56567 271
rect 56645 225 56691 271
rect 56769 225 56815 271
rect 56893 225 56939 271
rect 57017 225 57063 271
rect 57141 225 57187 271
rect 57265 225 57311 271
rect 57389 225 57435 271
rect 57513 225 57559 271
rect 57637 225 57683 271
rect 57761 225 57807 271
rect 57885 225 57931 271
rect 58009 225 58055 271
rect 58133 225 58179 271
rect 58257 225 58303 271
rect 58381 225 58427 271
rect 58505 225 58551 271
rect 58629 225 58675 271
rect 58753 225 58799 271
rect 58877 225 58923 271
rect 59001 225 59047 271
rect 59125 225 59171 271
rect 59249 225 59295 271
rect 59373 225 59419 271
rect 59497 225 59543 271
rect 59621 225 59667 271
rect 59745 225 59791 271
rect 59869 225 59915 271
rect 59993 225 60039 271
rect 60117 225 60163 271
rect 60241 225 60287 271
rect 60365 225 60411 271
rect 60489 225 60535 271
rect 60613 225 60659 271
rect 60737 225 60783 271
rect 60861 225 60907 271
rect 60985 225 61031 271
rect 61109 225 61155 271
rect 61233 225 61279 271
rect 61357 225 61403 271
rect 61481 225 61527 271
rect 61605 225 61651 271
rect 61729 225 61775 271
rect 61853 225 61899 271
rect 61977 225 62023 271
rect 62101 225 62147 271
rect 62225 225 62271 271
rect 62349 225 62395 271
rect 62473 225 62519 271
rect 62597 225 62643 271
rect 62721 225 62767 271
rect 62845 225 62891 271
rect 62969 225 63015 271
rect 63093 225 63139 271
rect 63217 225 63263 271
rect 63341 225 63387 271
rect 63465 225 63511 271
rect 63589 225 63635 271
rect 63713 225 63759 271
rect 63837 225 63883 271
rect 63961 225 64007 271
rect 64085 225 64131 271
rect 64209 225 64255 271
rect 64333 225 64379 271
rect 64457 225 64503 271
rect 64581 225 64627 271
rect 64705 225 64751 271
rect 64829 225 64875 271
rect 64953 225 64999 271
rect 65077 225 65123 271
rect 65201 225 65247 271
rect 65325 225 65371 271
rect 65449 225 65495 271
rect 65573 225 65619 271
rect 65697 225 65743 271
rect 65821 225 65867 271
rect 65945 225 65991 271
rect 66069 225 66115 271
rect 66193 225 66239 271
rect 66317 225 66363 271
rect 66441 225 66487 271
rect 66565 225 66611 271
rect 66689 225 66735 271
rect 66813 225 66859 271
rect 66937 225 66983 271
rect 67061 225 67107 271
rect 67185 225 67231 271
rect 67309 225 67355 271
rect 67433 225 67479 271
rect 67557 225 67603 271
rect 67681 225 67727 271
rect 67805 225 67851 271
rect 67929 225 67975 271
rect 68053 225 68099 271
rect 68177 225 68223 271
rect 68301 225 68347 271
rect 68425 225 68471 271
rect 68549 225 68595 271
rect 68673 225 68719 271
rect 68797 225 68843 271
rect 68921 225 68967 271
rect 69045 225 69091 271
rect 69169 225 69215 271
rect 69293 225 69339 271
rect 69417 225 69463 271
rect 69541 225 69587 271
rect 69665 225 69711 271
rect 69789 225 69835 271
rect 69913 225 69959 271
rect 70037 225 70083 271
rect 70161 225 70207 271
rect 70285 225 70331 271
rect 70409 225 70455 271
rect 70533 225 70579 271
rect 70657 225 70703 271
rect 70781 225 70827 271
rect 70905 225 70951 271
rect 71029 225 71075 271
rect 71153 225 71199 271
rect 71277 225 71323 271
rect 71401 225 71447 271
rect 71525 225 71571 271
rect 71649 225 71695 271
rect 71773 225 71819 271
rect 71897 225 71943 271
rect 72021 225 72067 271
rect 72145 225 72191 271
rect 72269 225 72315 271
rect 72393 225 72439 271
rect 72517 225 72563 271
rect 72641 225 72687 271
rect 72765 225 72811 271
rect 72889 225 72935 271
rect 73013 225 73059 271
rect 73137 225 73183 271
rect 73261 225 73307 271
rect 73385 225 73431 271
rect 73509 225 73555 271
rect 73633 225 73679 271
rect 73757 225 73803 271
rect 73881 225 73927 271
rect 74005 225 74051 271
rect 74129 225 74175 271
rect 74253 225 74299 271
rect 74377 225 74423 271
rect 74501 225 74547 271
rect 74625 225 74671 271
rect 74749 225 74795 271
rect 74873 225 74919 271
rect 74997 225 75043 271
rect 75121 225 75167 271
rect 75245 225 75291 271
rect 75369 225 75415 271
rect 75493 225 75539 271
rect 75617 225 75663 271
rect 75741 225 75787 271
rect 75865 225 75911 271
rect 75989 225 76035 271
rect 76113 225 76159 271
rect 76237 225 76283 271
rect 76361 225 76407 271
rect 76485 225 76531 271
rect 76609 225 76655 271
rect 76733 225 76779 271
rect 76857 225 76903 271
rect 76981 225 77027 271
rect 77105 225 77151 271
rect 77229 225 77275 271
rect 77353 225 77399 271
rect 77477 225 77523 271
rect 77601 225 77647 271
rect 77725 225 77771 271
rect 77849 225 77895 271
rect 77973 225 78019 271
rect 78097 225 78143 271
rect 78221 225 78267 271
rect 78345 225 78391 271
rect 78469 225 78515 271
rect 78593 225 78639 271
rect 78717 225 78763 271
rect 78841 225 78887 271
rect 78965 225 79011 271
rect 79089 225 79135 271
rect 79213 225 79259 271
rect 79337 225 79383 271
rect 79461 225 79507 271
rect 79585 225 79631 271
rect 79709 225 79755 271
rect 79833 225 79879 271
rect 79957 225 80003 271
rect 80081 225 80127 271
rect 80205 225 80251 271
rect 80329 225 80375 271
rect 80453 225 80499 271
rect 80577 225 80623 271
rect 80701 225 80747 271
rect 80825 225 80871 271
rect 80949 225 80995 271
rect 81073 225 81119 271
rect 81197 225 81243 271
rect 81321 225 81367 271
rect 81445 225 81491 271
rect 81569 225 81615 271
rect 81693 225 81739 271
rect 81817 225 81863 271
rect 81941 225 81987 271
rect 82065 225 82111 271
rect 82189 225 82235 271
rect 82313 225 82359 271
rect 82437 225 82483 271
rect 82561 225 82607 271
rect 82685 225 82731 271
rect 82809 225 82855 271
rect 82933 225 82979 271
rect 83057 225 83103 271
rect 83181 225 83227 271
rect 83305 225 83351 271
rect 83429 225 83475 271
rect 83553 225 83599 271
rect 83677 225 83723 271
rect 83801 225 83847 271
rect 83925 225 83971 271
rect 84049 225 84095 271
rect 84173 225 84219 271
rect 84297 225 84343 271
rect 84421 225 84467 271
rect 84545 225 84591 271
rect 84669 225 84715 271
rect 84793 225 84839 271
rect 84917 225 84963 271
rect 85041 225 85087 271
rect 85165 225 85211 271
rect 85289 225 85335 271
rect 85413 225 85459 271
rect 85537 225 85583 271
rect -23 101 23 147
rect 101 101 147 147
rect 225 101 271 147
rect 349 101 395 147
rect 473 101 519 147
rect 597 101 643 147
rect 721 101 767 147
rect 845 101 891 147
rect 969 101 1015 147
rect 1093 101 1139 147
rect 1217 101 1263 147
rect 1341 101 1387 147
rect 1465 101 1511 147
rect 1589 101 1635 147
rect 1713 101 1759 147
rect 1837 101 1883 147
rect 1961 101 2007 147
rect 2085 101 2131 147
rect 2209 101 2255 147
rect 2333 101 2379 147
rect 2457 101 2503 147
rect 2581 101 2627 147
rect 2705 101 2751 147
rect 2829 101 2875 147
rect 2953 101 2999 147
rect 3077 101 3123 147
rect 3201 101 3247 147
rect 3325 101 3371 147
rect 3449 101 3495 147
rect 3573 101 3619 147
rect 3697 101 3743 147
rect 3821 101 3867 147
rect 3945 101 3991 147
rect 4069 101 4115 147
rect 4193 101 4239 147
rect 4317 101 4363 147
rect 4441 101 4487 147
rect 4565 101 4611 147
rect 4689 101 4735 147
rect 4813 101 4859 147
rect 4937 101 4983 147
rect 5061 101 5107 147
rect 5185 101 5231 147
rect 5309 101 5355 147
rect 5433 101 5479 147
rect 5557 101 5603 147
rect 5681 101 5727 147
rect 5805 101 5851 147
rect 5929 101 5975 147
rect 6053 101 6099 147
rect 6177 101 6223 147
rect 6301 101 6347 147
rect 6425 101 6471 147
rect 6549 101 6595 147
rect 6673 101 6719 147
rect 6797 101 6843 147
rect 6921 101 6967 147
rect 7045 101 7091 147
rect 7169 101 7215 147
rect 7293 101 7339 147
rect 7417 101 7463 147
rect 7541 101 7587 147
rect 7665 101 7711 147
rect 7789 101 7835 147
rect 7913 101 7959 147
rect 8037 101 8083 147
rect 8161 101 8207 147
rect 8285 101 8331 147
rect 8409 101 8455 147
rect 8533 101 8579 147
rect 8657 101 8703 147
rect 8781 101 8827 147
rect 8905 101 8951 147
rect 9029 101 9075 147
rect 9153 101 9199 147
rect 9277 101 9323 147
rect 9401 101 9447 147
rect 9525 101 9571 147
rect 9649 101 9695 147
rect 9773 101 9819 147
rect 9897 101 9943 147
rect 10021 101 10067 147
rect 10145 101 10191 147
rect 10269 101 10315 147
rect 10393 101 10439 147
rect 10517 101 10563 147
rect 10641 101 10687 147
rect 10765 101 10811 147
rect 10889 101 10935 147
rect 11013 101 11059 147
rect 11137 101 11183 147
rect 11261 101 11307 147
rect 11385 101 11431 147
rect 11509 101 11555 147
rect 11633 101 11679 147
rect 11757 101 11803 147
rect 11881 101 11927 147
rect 12005 101 12051 147
rect 12129 101 12175 147
rect 12253 101 12299 147
rect 12377 101 12423 147
rect 12501 101 12547 147
rect 12625 101 12671 147
rect 12749 101 12795 147
rect 12873 101 12919 147
rect 12997 101 13043 147
rect 13121 101 13167 147
rect 13245 101 13291 147
rect 13369 101 13415 147
rect 13493 101 13539 147
rect 13617 101 13663 147
rect 13741 101 13787 147
rect 13865 101 13911 147
rect 13989 101 14035 147
rect 14113 101 14159 147
rect 14237 101 14283 147
rect 14361 101 14407 147
rect 14485 101 14531 147
rect 14609 101 14655 147
rect 14733 101 14779 147
rect 14857 101 14903 147
rect 14981 101 15027 147
rect 15105 101 15151 147
rect 15229 101 15275 147
rect 15353 101 15399 147
rect 15477 101 15523 147
rect 15601 101 15647 147
rect 15725 101 15771 147
rect 15849 101 15895 147
rect 15973 101 16019 147
rect 16097 101 16143 147
rect 16221 101 16267 147
rect 16345 101 16391 147
rect 16469 101 16515 147
rect 16593 101 16639 147
rect 16717 101 16763 147
rect 16841 101 16887 147
rect 16965 101 17011 147
rect 17089 101 17135 147
rect 17213 101 17259 147
rect 17337 101 17383 147
rect 17461 101 17507 147
rect 17585 101 17631 147
rect 17709 101 17755 147
rect 17833 101 17879 147
rect 17957 101 18003 147
rect 18081 101 18127 147
rect 18205 101 18251 147
rect 18329 101 18375 147
rect 18453 101 18499 147
rect 18577 101 18623 147
rect 18701 101 18747 147
rect 18825 101 18871 147
rect 18949 101 18995 147
rect 19073 101 19119 147
rect 19197 101 19243 147
rect 19321 101 19367 147
rect 19445 101 19491 147
rect 19569 101 19615 147
rect 19693 101 19739 147
rect 19817 101 19863 147
rect 19941 101 19987 147
rect 20065 101 20111 147
rect 20189 101 20235 147
rect 20313 101 20359 147
rect 20437 101 20483 147
rect 20561 101 20607 147
rect 20685 101 20731 147
rect 20809 101 20855 147
rect 20933 101 20979 147
rect 21057 101 21103 147
rect 21181 101 21227 147
rect 21305 101 21351 147
rect 21429 101 21475 147
rect 21553 101 21599 147
rect 21677 101 21723 147
rect 21801 101 21847 147
rect 21925 101 21971 147
rect 22049 101 22095 147
rect 22173 101 22219 147
rect 22297 101 22343 147
rect 22421 101 22467 147
rect 22545 101 22591 147
rect 22669 101 22715 147
rect 22793 101 22839 147
rect 22917 101 22963 147
rect 23041 101 23087 147
rect 23165 101 23211 147
rect 23289 101 23335 147
rect 23413 101 23459 147
rect 23537 101 23583 147
rect 23661 101 23707 147
rect 23785 101 23831 147
rect 23909 101 23955 147
rect 24033 101 24079 147
rect 24157 101 24203 147
rect 24281 101 24327 147
rect 24405 101 24451 147
rect 24529 101 24575 147
rect 24653 101 24699 147
rect 24777 101 24823 147
rect 24901 101 24947 147
rect 25025 101 25071 147
rect 25149 101 25195 147
rect 25273 101 25319 147
rect 25397 101 25443 147
rect 25521 101 25567 147
rect 25645 101 25691 147
rect 25769 101 25815 147
rect 25893 101 25939 147
rect 26017 101 26063 147
rect 26141 101 26187 147
rect 26265 101 26311 147
rect 26389 101 26435 147
rect 26513 101 26559 147
rect 26637 101 26683 147
rect 26761 101 26807 147
rect 26885 101 26931 147
rect 27009 101 27055 147
rect 27133 101 27179 147
rect 27257 101 27303 147
rect 27381 101 27427 147
rect 27505 101 27551 147
rect 27629 101 27675 147
rect 27753 101 27799 147
rect 27877 101 27923 147
rect 28001 101 28047 147
rect 28125 101 28171 147
rect 28249 101 28295 147
rect 28373 101 28419 147
rect 28497 101 28543 147
rect 28621 101 28667 147
rect 28745 101 28791 147
rect 28869 101 28915 147
rect 28993 101 29039 147
rect 29117 101 29163 147
rect 29241 101 29287 147
rect 29365 101 29411 147
rect 29489 101 29535 147
rect 29613 101 29659 147
rect 29737 101 29783 147
rect 29861 101 29907 147
rect 29985 101 30031 147
rect 30109 101 30155 147
rect 30233 101 30279 147
rect 30357 101 30403 147
rect 30481 101 30527 147
rect 30605 101 30651 147
rect 30729 101 30775 147
rect 30853 101 30899 147
rect 30977 101 31023 147
rect 31101 101 31147 147
rect 31225 101 31271 147
rect 31349 101 31395 147
rect 31473 101 31519 147
rect 31597 101 31643 147
rect 31721 101 31767 147
rect 31845 101 31891 147
rect 31969 101 32015 147
rect 32093 101 32139 147
rect 32217 101 32263 147
rect 32341 101 32387 147
rect 32465 101 32511 147
rect 32589 101 32635 147
rect 32713 101 32759 147
rect 32837 101 32883 147
rect 32961 101 33007 147
rect 33085 101 33131 147
rect 33209 101 33255 147
rect 33333 101 33379 147
rect 33457 101 33503 147
rect 33581 101 33627 147
rect 33705 101 33751 147
rect 33829 101 33875 147
rect 33953 101 33999 147
rect 34077 101 34123 147
rect 34201 101 34247 147
rect 34325 101 34371 147
rect 34449 101 34495 147
rect 34573 101 34619 147
rect 34697 101 34743 147
rect 34821 101 34867 147
rect 34945 101 34991 147
rect 35069 101 35115 147
rect 35193 101 35239 147
rect 35317 101 35363 147
rect 35441 101 35487 147
rect 35565 101 35611 147
rect 35689 101 35735 147
rect 35813 101 35859 147
rect 35937 101 35983 147
rect 36061 101 36107 147
rect 36185 101 36231 147
rect 36309 101 36355 147
rect 36433 101 36479 147
rect 36557 101 36603 147
rect 36681 101 36727 147
rect 36805 101 36851 147
rect 36929 101 36975 147
rect 37053 101 37099 147
rect 37177 101 37223 147
rect 37301 101 37347 147
rect 37425 101 37471 147
rect 37549 101 37595 147
rect 37673 101 37719 147
rect 37797 101 37843 147
rect 37921 101 37967 147
rect 38045 101 38091 147
rect 38169 101 38215 147
rect 38293 101 38339 147
rect 38417 101 38463 147
rect 38541 101 38587 147
rect 38665 101 38711 147
rect 38789 101 38835 147
rect 38913 101 38959 147
rect 39037 101 39083 147
rect 39161 101 39207 147
rect 39285 101 39331 147
rect 39409 101 39455 147
rect 39533 101 39579 147
rect 39657 101 39703 147
rect 39781 101 39827 147
rect 39905 101 39951 147
rect 40029 101 40075 147
rect 40153 101 40199 147
rect 40277 101 40323 147
rect 40401 101 40447 147
rect 40525 101 40571 147
rect 40649 101 40695 147
rect 40773 101 40819 147
rect 40897 101 40943 147
rect 41021 101 41067 147
rect 41145 101 41191 147
rect 41269 101 41315 147
rect 41393 101 41439 147
rect 41517 101 41563 147
rect 41641 101 41687 147
rect 41765 101 41811 147
rect 41889 101 41935 147
rect 42013 101 42059 147
rect 42137 101 42183 147
rect 42261 101 42307 147
rect 42385 101 42431 147
rect 42509 101 42555 147
rect 42633 101 42679 147
rect 42757 101 42803 147
rect 42881 101 42927 147
rect 43005 101 43051 147
rect 43129 101 43175 147
rect 43253 101 43299 147
rect 43377 101 43423 147
rect 43501 101 43547 147
rect 43625 101 43671 147
rect 43749 101 43795 147
rect 43873 101 43919 147
rect 43997 101 44043 147
rect 44121 101 44167 147
rect 44245 101 44291 147
rect 44369 101 44415 147
rect 44493 101 44539 147
rect 44617 101 44663 147
rect 44741 101 44787 147
rect 44865 101 44911 147
rect 44989 101 45035 147
rect 45113 101 45159 147
rect 45237 101 45283 147
rect 45361 101 45407 147
rect 45485 101 45531 147
rect 45609 101 45655 147
rect 45733 101 45779 147
rect 45857 101 45903 147
rect 45981 101 46027 147
rect 46105 101 46151 147
rect 46229 101 46275 147
rect 46353 101 46399 147
rect 46477 101 46523 147
rect 46601 101 46647 147
rect 46725 101 46771 147
rect 46849 101 46895 147
rect 46973 101 47019 147
rect 47097 101 47143 147
rect 47221 101 47267 147
rect 47345 101 47391 147
rect 47469 101 47515 147
rect 47593 101 47639 147
rect 47717 101 47763 147
rect 47841 101 47887 147
rect 47965 101 48011 147
rect 48089 101 48135 147
rect 48213 101 48259 147
rect 48337 101 48383 147
rect 48461 101 48507 147
rect 48585 101 48631 147
rect 48709 101 48755 147
rect 48833 101 48879 147
rect 48957 101 49003 147
rect 49081 101 49127 147
rect 49205 101 49251 147
rect 49329 101 49375 147
rect 49453 101 49499 147
rect 49577 101 49623 147
rect 49701 101 49747 147
rect 49825 101 49871 147
rect 49949 101 49995 147
rect 50073 101 50119 147
rect 50197 101 50243 147
rect 50321 101 50367 147
rect 50445 101 50491 147
rect 50569 101 50615 147
rect 50693 101 50739 147
rect 50817 101 50863 147
rect 50941 101 50987 147
rect 51065 101 51111 147
rect 51189 101 51235 147
rect 51313 101 51359 147
rect 51437 101 51483 147
rect 51561 101 51607 147
rect 51685 101 51731 147
rect 51809 101 51855 147
rect 51933 101 51979 147
rect 52057 101 52103 147
rect 52181 101 52227 147
rect 52305 101 52351 147
rect 52429 101 52475 147
rect 52553 101 52599 147
rect 52677 101 52723 147
rect 52801 101 52847 147
rect 52925 101 52971 147
rect 53049 101 53095 147
rect 53173 101 53219 147
rect 53297 101 53343 147
rect 53421 101 53467 147
rect 53545 101 53591 147
rect 53669 101 53715 147
rect 53793 101 53839 147
rect 53917 101 53963 147
rect 54041 101 54087 147
rect 54165 101 54211 147
rect 54289 101 54335 147
rect 54413 101 54459 147
rect 54537 101 54583 147
rect 54661 101 54707 147
rect 54785 101 54831 147
rect 54909 101 54955 147
rect 55033 101 55079 147
rect 55157 101 55203 147
rect 55281 101 55327 147
rect 55405 101 55451 147
rect 55529 101 55575 147
rect 55653 101 55699 147
rect 55777 101 55823 147
rect 55901 101 55947 147
rect 56025 101 56071 147
rect 56149 101 56195 147
rect 56273 101 56319 147
rect 56397 101 56443 147
rect 56521 101 56567 147
rect 56645 101 56691 147
rect 56769 101 56815 147
rect 56893 101 56939 147
rect 57017 101 57063 147
rect 57141 101 57187 147
rect 57265 101 57311 147
rect 57389 101 57435 147
rect 57513 101 57559 147
rect 57637 101 57683 147
rect 57761 101 57807 147
rect 57885 101 57931 147
rect 58009 101 58055 147
rect 58133 101 58179 147
rect 58257 101 58303 147
rect 58381 101 58427 147
rect 58505 101 58551 147
rect 58629 101 58675 147
rect 58753 101 58799 147
rect 58877 101 58923 147
rect 59001 101 59047 147
rect 59125 101 59171 147
rect 59249 101 59295 147
rect 59373 101 59419 147
rect 59497 101 59543 147
rect 59621 101 59667 147
rect 59745 101 59791 147
rect 59869 101 59915 147
rect 59993 101 60039 147
rect 60117 101 60163 147
rect 60241 101 60287 147
rect 60365 101 60411 147
rect 60489 101 60535 147
rect 60613 101 60659 147
rect 60737 101 60783 147
rect 60861 101 60907 147
rect 60985 101 61031 147
rect 61109 101 61155 147
rect 61233 101 61279 147
rect 61357 101 61403 147
rect 61481 101 61527 147
rect 61605 101 61651 147
rect 61729 101 61775 147
rect 61853 101 61899 147
rect 61977 101 62023 147
rect 62101 101 62147 147
rect 62225 101 62271 147
rect 62349 101 62395 147
rect 62473 101 62519 147
rect 62597 101 62643 147
rect 62721 101 62767 147
rect 62845 101 62891 147
rect 62969 101 63015 147
rect 63093 101 63139 147
rect 63217 101 63263 147
rect 63341 101 63387 147
rect 63465 101 63511 147
rect 63589 101 63635 147
rect 63713 101 63759 147
rect 63837 101 63883 147
rect 63961 101 64007 147
rect 64085 101 64131 147
rect 64209 101 64255 147
rect 64333 101 64379 147
rect 64457 101 64503 147
rect 64581 101 64627 147
rect 64705 101 64751 147
rect 64829 101 64875 147
rect 64953 101 64999 147
rect 65077 101 65123 147
rect 65201 101 65247 147
rect 65325 101 65371 147
rect 65449 101 65495 147
rect 65573 101 65619 147
rect 65697 101 65743 147
rect 65821 101 65867 147
rect 65945 101 65991 147
rect 66069 101 66115 147
rect 66193 101 66239 147
rect 66317 101 66363 147
rect 66441 101 66487 147
rect 66565 101 66611 147
rect 66689 101 66735 147
rect 66813 101 66859 147
rect 66937 101 66983 147
rect 67061 101 67107 147
rect 67185 101 67231 147
rect 67309 101 67355 147
rect 67433 101 67479 147
rect 67557 101 67603 147
rect 67681 101 67727 147
rect 67805 101 67851 147
rect 67929 101 67975 147
rect 68053 101 68099 147
rect 68177 101 68223 147
rect 68301 101 68347 147
rect 68425 101 68471 147
rect 68549 101 68595 147
rect 68673 101 68719 147
rect 68797 101 68843 147
rect 68921 101 68967 147
rect 69045 101 69091 147
rect 69169 101 69215 147
rect 69293 101 69339 147
rect 69417 101 69463 147
rect 69541 101 69587 147
rect 69665 101 69711 147
rect 69789 101 69835 147
rect 69913 101 69959 147
rect 70037 101 70083 147
rect 70161 101 70207 147
rect 70285 101 70331 147
rect 70409 101 70455 147
rect 70533 101 70579 147
rect 70657 101 70703 147
rect 70781 101 70827 147
rect 70905 101 70951 147
rect 71029 101 71075 147
rect 71153 101 71199 147
rect 71277 101 71323 147
rect 71401 101 71447 147
rect 71525 101 71571 147
rect 71649 101 71695 147
rect 71773 101 71819 147
rect 71897 101 71943 147
rect 72021 101 72067 147
rect 72145 101 72191 147
rect 72269 101 72315 147
rect 72393 101 72439 147
rect 72517 101 72563 147
rect 72641 101 72687 147
rect 72765 101 72811 147
rect 72889 101 72935 147
rect 73013 101 73059 147
rect 73137 101 73183 147
rect 73261 101 73307 147
rect 73385 101 73431 147
rect 73509 101 73555 147
rect 73633 101 73679 147
rect 73757 101 73803 147
rect 73881 101 73927 147
rect 74005 101 74051 147
rect 74129 101 74175 147
rect 74253 101 74299 147
rect 74377 101 74423 147
rect 74501 101 74547 147
rect 74625 101 74671 147
rect 74749 101 74795 147
rect 74873 101 74919 147
rect 74997 101 75043 147
rect 75121 101 75167 147
rect 75245 101 75291 147
rect 75369 101 75415 147
rect 75493 101 75539 147
rect 75617 101 75663 147
rect 75741 101 75787 147
rect 75865 101 75911 147
rect 75989 101 76035 147
rect 76113 101 76159 147
rect 76237 101 76283 147
rect 76361 101 76407 147
rect 76485 101 76531 147
rect 76609 101 76655 147
rect 76733 101 76779 147
rect 76857 101 76903 147
rect 76981 101 77027 147
rect 77105 101 77151 147
rect 77229 101 77275 147
rect 77353 101 77399 147
rect 77477 101 77523 147
rect 77601 101 77647 147
rect 77725 101 77771 147
rect 77849 101 77895 147
rect 77973 101 78019 147
rect 78097 101 78143 147
rect 78221 101 78267 147
rect 78345 101 78391 147
rect 78469 101 78515 147
rect 78593 101 78639 147
rect 78717 101 78763 147
rect 78841 101 78887 147
rect 78965 101 79011 147
rect 79089 101 79135 147
rect 79213 101 79259 147
rect 79337 101 79383 147
rect 79461 101 79507 147
rect 79585 101 79631 147
rect 79709 101 79755 147
rect 79833 101 79879 147
rect 79957 101 80003 147
rect 80081 101 80127 147
rect 80205 101 80251 147
rect 80329 101 80375 147
rect 80453 101 80499 147
rect 80577 101 80623 147
rect 80701 101 80747 147
rect 80825 101 80871 147
rect 80949 101 80995 147
rect 81073 101 81119 147
rect 81197 101 81243 147
rect 81321 101 81367 147
rect 81445 101 81491 147
rect 81569 101 81615 147
rect 81693 101 81739 147
rect 81817 101 81863 147
rect 81941 101 81987 147
rect 82065 101 82111 147
rect 82189 101 82235 147
rect 82313 101 82359 147
rect 82437 101 82483 147
rect 82561 101 82607 147
rect 82685 101 82731 147
rect 82809 101 82855 147
rect 82933 101 82979 147
rect 83057 101 83103 147
rect 83181 101 83227 147
rect 83305 101 83351 147
rect 83429 101 83475 147
rect 83553 101 83599 147
rect 83677 101 83723 147
rect 83801 101 83847 147
rect 83925 101 83971 147
rect 84049 101 84095 147
rect 84173 101 84219 147
rect 84297 101 84343 147
rect 84421 101 84467 147
rect 84545 101 84591 147
rect 84669 101 84715 147
rect 84793 101 84839 147
rect 84917 101 84963 147
rect 85041 101 85087 147
rect 85165 101 85211 147
rect 85289 101 85335 147
rect 85413 101 85459 147
rect 85537 101 85583 147
rect -23 -23 23 23
rect 101 -23 147 23
rect 225 -23 271 23
rect 349 -23 395 23
rect 473 -23 519 23
rect 597 -23 643 23
rect 721 -23 767 23
rect 845 -23 891 23
rect 969 -23 1015 23
rect 1093 -23 1139 23
rect 1217 -23 1263 23
rect 1341 -23 1387 23
rect 1465 -23 1511 23
rect 1589 -23 1635 23
rect 1713 -23 1759 23
rect 1837 -23 1883 23
rect 1961 -23 2007 23
rect 2085 -23 2131 23
rect 2209 -23 2255 23
rect 2333 -23 2379 23
rect 2457 -23 2503 23
rect 2581 -23 2627 23
rect 2705 -23 2751 23
rect 2829 -23 2875 23
rect 2953 -23 2999 23
rect 3077 -23 3123 23
rect 3201 -23 3247 23
rect 3325 -23 3371 23
rect 3449 -23 3495 23
rect 3573 -23 3619 23
rect 3697 -23 3743 23
rect 3821 -23 3867 23
rect 3945 -23 3991 23
rect 4069 -23 4115 23
rect 4193 -23 4239 23
rect 4317 -23 4363 23
rect 4441 -23 4487 23
rect 4565 -23 4611 23
rect 4689 -23 4735 23
rect 4813 -23 4859 23
rect 4937 -23 4983 23
rect 5061 -23 5107 23
rect 5185 -23 5231 23
rect 5309 -23 5355 23
rect 5433 -23 5479 23
rect 5557 -23 5603 23
rect 5681 -23 5727 23
rect 5805 -23 5851 23
rect 5929 -23 5975 23
rect 6053 -23 6099 23
rect 6177 -23 6223 23
rect 6301 -23 6347 23
rect 6425 -23 6471 23
rect 6549 -23 6595 23
rect 6673 -23 6719 23
rect 6797 -23 6843 23
rect 6921 -23 6967 23
rect 7045 -23 7091 23
rect 7169 -23 7215 23
rect 7293 -23 7339 23
rect 7417 -23 7463 23
rect 7541 -23 7587 23
rect 7665 -23 7711 23
rect 7789 -23 7835 23
rect 7913 -23 7959 23
rect 8037 -23 8083 23
rect 8161 -23 8207 23
rect 8285 -23 8331 23
rect 8409 -23 8455 23
rect 8533 -23 8579 23
rect 8657 -23 8703 23
rect 8781 -23 8827 23
rect 8905 -23 8951 23
rect 9029 -23 9075 23
rect 9153 -23 9199 23
rect 9277 -23 9323 23
rect 9401 -23 9447 23
rect 9525 -23 9571 23
rect 9649 -23 9695 23
rect 9773 -23 9819 23
rect 9897 -23 9943 23
rect 10021 -23 10067 23
rect 10145 -23 10191 23
rect 10269 -23 10315 23
rect 10393 -23 10439 23
rect 10517 -23 10563 23
rect 10641 -23 10687 23
rect 10765 -23 10811 23
rect 10889 -23 10935 23
rect 11013 -23 11059 23
rect 11137 -23 11183 23
rect 11261 -23 11307 23
rect 11385 -23 11431 23
rect 11509 -23 11555 23
rect 11633 -23 11679 23
rect 11757 -23 11803 23
rect 11881 -23 11927 23
rect 12005 -23 12051 23
rect 12129 -23 12175 23
rect 12253 -23 12299 23
rect 12377 -23 12423 23
rect 12501 -23 12547 23
rect 12625 -23 12671 23
rect 12749 -23 12795 23
rect 12873 -23 12919 23
rect 12997 -23 13043 23
rect 13121 -23 13167 23
rect 13245 -23 13291 23
rect 13369 -23 13415 23
rect 13493 -23 13539 23
rect 13617 -23 13663 23
rect 13741 -23 13787 23
rect 13865 -23 13911 23
rect 13989 -23 14035 23
rect 14113 -23 14159 23
rect 14237 -23 14283 23
rect 14361 -23 14407 23
rect 14485 -23 14531 23
rect 14609 -23 14655 23
rect 14733 -23 14779 23
rect 14857 -23 14903 23
rect 14981 -23 15027 23
rect 15105 -23 15151 23
rect 15229 -23 15275 23
rect 15353 -23 15399 23
rect 15477 -23 15523 23
rect 15601 -23 15647 23
rect 15725 -23 15771 23
rect 15849 -23 15895 23
rect 15973 -23 16019 23
rect 16097 -23 16143 23
rect 16221 -23 16267 23
rect 16345 -23 16391 23
rect 16469 -23 16515 23
rect 16593 -23 16639 23
rect 16717 -23 16763 23
rect 16841 -23 16887 23
rect 16965 -23 17011 23
rect 17089 -23 17135 23
rect 17213 -23 17259 23
rect 17337 -23 17383 23
rect 17461 -23 17507 23
rect 17585 -23 17631 23
rect 17709 -23 17755 23
rect 17833 -23 17879 23
rect 17957 -23 18003 23
rect 18081 -23 18127 23
rect 18205 -23 18251 23
rect 18329 -23 18375 23
rect 18453 -23 18499 23
rect 18577 -23 18623 23
rect 18701 -23 18747 23
rect 18825 -23 18871 23
rect 18949 -23 18995 23
rect 19073 -23 19119 23
rect 19197 -23 19243 23
rect 19321 -23 19367 23
rect 19445 -23 19491 23
rect 19569 -23 19615 23
rect 19693 -23 19739 23
rect 19817 -23 19863 23
rect 19941 -23 19987 23
rect 20065 -23 20111 23
rect 20189 -23 20235 23
rect 20313 -23 20359 23
rect 20437 -23 20483 23
rect 20561 -23 20607 23
rect 20685 -23 20731 23
rect 20809 -23 20855 23
rect 20933 -23 20979 23
rect 21057 -23 21103 23
rect 21181 -23 21227 23
rect 21305 -23 21351 23
rect 21429 -23 21475 23
rect 21553 -23 21599 23
rect 21677 -23 21723 23
rect 21801 -23 21847 23
rect 21925 -23 21971 23
rect 22049 -23 22095 23
rect 22173 -23 22219 23
rect 22297 -23 22343 23
rect 22421 -23 22467 23
rect 22545 -23 22591 23
rect 22669 -23 22715 23
rect 22793 -23 22839 23
rect 22917 -23 22963 23
rect 23041 -23 23087 23
rect 23165 -23 23211 23
rect 23289 -23 23335 23
rect 23413 -23 23459 23
rect 23537 -23 23583 23
rect 23661 -23 23707 23
rect 23785 -23 23831 23
rect 23909 -23 23955 23
rect 24033 -23 24079 23
rect 24157 -23 24203 23
rect 24281 -23 24327 23
rect 24405 -23 24451 23
rect 24529 -23 24575 23
rect 24653 -23 24699 23
rect 24777 -23 24823 23
rect 24901 -23 24947 23
rect 25025 -23 25071 23
rect 25149 -23 25195 23
rect 25273 -23 25319 23
rect 25397 -23 25443 23
rect 25521 -23 25567 23
rect 25645 -23 25691 23
rect 25769 -23 25815 23
rect 25893 -23 25939 23
rect 26017 -23 26063 23
rect 26141 -23 26187 23
rect 26265 -23 26311 23
rect 26389 -23 26435 23
rect 26513 -23 26559 23
rect 26637 -23 26683 23
rect 26761 -23 26807 23
rect 26885 -23 26931 23
rect 27009 -23 27055 23
rect 27133 -23 27179 23
rect 27257 -23 27303 23
rect 27381 -23 27427 23
rect 27505 -23 27551 23
rect 27629 -23 27675 23
rect 27753 -23 27799 23
rect 27877 -23 27923 23
rect 28001 -23 28047 23
rect 28125 -23 28171 23
rect 28249 -23 28295 23
rect 28373 -23 28419 23
rect 28497 -23 28543 23
rect 28621 -23 28667 23
rect 28745 -23 28791 23
rect 28869 -23 28915 23
rect 28993 -23 29039 23
rect 29117 -23 29163 23
rect 29241 -23 29287 23
rect 29365 -23 29411 23
rect 29489 -23 29535 23
rect 29613 -23 29659 23
rect 29737 -23 29783 23
rect 29861 -23 29907 23
rect 29985 -23 30031 23
rect 30109 -23 30155 23
rect 30233 -23 30279 23
rect 30357 -23 30403 23
rect 30481 -23 30527 23
rect 30605 -23 30651 23
rect 30729 -23 30775 23
rect 30853 -23 30899 23
rect 30977 -23 31023 23
rect 31101 -23 31147 23
rect 31225 -23 31271 23
rect 31349 -23 31395 23
rect 31473 -23 31519 23
rect 31597 -23 31643 23
rect 31721 -23 31767 23
rect 31845 -23 31891 23
rect 31969 -23 32015 23
rect 32093 -23 32139 23
rect 32217 -23 32263 23
rect 32341 -23 32387 23
rect 32465 -23 32511 23
rect 32589 -23 32635 23
rect 32713 -23 32759 23
rect 32837 -23 32883 23
rect 32961 -23 33007 23
rect 33085 -23 33131 23
rect 33209 -23 33255 23
rect 33333 -23 33379 23
rect 33457 -23 33503 23
rect 33581 -23 33627 23
rect 33705 -23 33751 23
rect 33829 -23 33875 23
rect 33953 -23 33999 23
rect 34077 -23 34123 23
rect 34201 -23 34247 23
rect 34325 -23 34371 23
rect 34449 -23 34495 23
rect 34573 -23 34619 23
rect 34697 -23 34743 23
rect 34821 -23 34867 23
rect 34945 -23 34991 23
rect 35069 -23 35115 23
rect 35193 -23 35239 23
rect 35317 -23 35363 23
rect 35441 -23 35487 23
rect 35565 -23 35611 23
rect 35689 -23 35735 23
rect 35813 -23 35859 23
rect 35937 -23 35983 23
rect 36061 -23 36107 23
rect 36185 -23 36231 23
rect 36309 -23 36355 23
rect 36433 -23 36479 23
rect 36557 -23 36603 23
rect 36681 -23 36727 23
rect 36805 -23 36851 23
rect 36929 -23 36975 23
rect 37053 -23 37099 23
rect 37177 -23 37223 23
rect 37301 -23 37347 23
rect 37425 -23 37471 23
rect 37549 -23 37595 23
rect 37673 -23 37719 23
rect 37797 -23 37843 23
rect 37921 -23 37967 23
rect 38045 -23 38091 23
rect 38169 -23 38215 23
rect 38293 -23 38339 23
rect 38417 -23 38463 23
rect 38541 -23 38587 23
rect 38665 -23 38711 23
rect 38789 -23 38835 23
rect 38913 -23 38959 23
rect 39037 -23 39083 23
rect 39161 -23 39207 23
rect 39285 -23 39331 23
rect 39409 -23 39455 23
rect 39533 -23 39579 23
rect 39657 -23 39703 23
rect 39781 -23 39827 23
rect 39905 -23 39951 23
rect 40029 -23 40075 23
rect 40153 -23 40199 23
rect 40277 -23 40323 23
rect 40401 -23 40447 23
rect 40525 -23 40571 23
rect 40649 -23 40695 23
rect 40773 -23 40819 23
rect 40897 -23 40943 23
rect 41021 -23 41067 23
rect 41145 -23 41191 23
rect 41269 -23 41315 23
rect 41393 -23 41439 23
rect 41517 -23 41563 23
rect 41641 -23 41687 23
rect 41765 -23 41811 23
rect 41889 -23 41935 23
rect 42013 -23 42059 23
rect 42137 -23 42183 23
rect 42261 -23 42307 23
rect 42385 -23 42431 23
rect 42509 -23 42555 23
rect 42633 -23 42679 23
rect 42757 -23 42803 23
rect 42881 -23 42927 23
rect 43005 -23 43051 23
rect 43129 -23 43175 23
rect 43253 -23 43299 23
rect 43377 -23 43423 23
rect 43501 -23 43547 23
rect 43625 -23 43671 23
rect 43749 -23 43795 23
rect 43873 -23 43919 23
rect 43997 -23 44043 23
rect 44121 -23 44167 23
rect 44245 -23 44291 23
rect 44369 -23 44415 23
rect 44493 -23 44539 23
rect 44617 -23 44663 23
rect 44741 -23 44787 23
rect 44865 -23 44911 23
rect 44989 -23 45035 23
rect 45113 -23 45159 23
rect 45237 -23 45283 23
rect 45361 -23 45407 23
rect 45485 -23 45531 23
rect 45609 -23 45655 23
rect 45733 -23 45779 23
rect 45857 -23 45903 23
rect 45981 -23 46027 23
rect 46105 -23 46151 23
rect 46229 -23 46275 23
rect 46353 -23 46399 23
rect 46477 -23 46523 23
rect 46601 -23 46647 23
rect 46725 -23 46771 23
rect 46849 -23 46895 23
rect 46973 -23 47019 23
rect 47097 -23 47143 23
rect 47221 -23 47267 23
rect 47345 -23 47391 23
rect 47469 -23 47515 23
rect 47593 -23 47639 23
rect 47717 -23 47763 23
rect 47841 -23 47887 23
rect 47965 -23 48011 23
rect 48089 -23 48135 23
rect 48213 -23 48259 23
rect 48337 -23 48383 23
rect 48461 -23 48507 23
rect 48585 -23 48631 23
rect 48709 -23 48755 23
rect 48833 -23 48879 23
rect 48957 -23 49003 23
rect 49081 -23 49127 23
rect 49205 -23 49251 23
rect 49329 -23 49375 23
rect 49453 -23 49499 23
rect 49577 -23 49623 23
rect 49701 -23 49747 23
rect 49825 -23 49871 23
rect 49949 -23 49995 23
rect 50073 -23 50119 23
rect 50197 -23 50243 23
rect 50321 -23 50367 23
rect 50445 -23 50491 23
rect 50569 -23 50615 23
rect 50693 -23 50739 23
rect 50817 -23 50863 23
rect 50941 -23 50987 23
rect 51065 -23 51111 23
rect 51189 -23 51235 23
rect 51313 -23 51359 23
rect 51437 -23 51483 23
rect 51561 -23 51607 23
rect 51685 -23 51731 23
rect 51809 -23 51855 23
rect 51933 -23 51979 23
rect 52057 -23 52103 23
rect 52181 -23 52227 23
rect 52305 -23 52351 23
rect 52429 -23 52475 23
rect 52553 -23 52599 23
rect 52677 -23 52723 23
rect 52801 -23 52847 23
rect 52925 -23 52971 23
rect 53049 -23 53095 23
rect 53173 -23 53219 23
rect 53297 -23 53343 23
rect 53421 -23 53467 23
rect 53545 -23 53591 23
rect 53669 -23 53715 23
rect 53793 -23 53839 23
rect 53917 -23 53963 23
rect 54041 -23 54087 23
rect 54165 -23 54211 23
rect 54289 -23 54335 23
rect 54413 -23 54459 23
rect 54537 -23 54583 23
rect 54661 -23 54707 23
rect 54785 -23 54831 23
rect 54909 -23 54955 23
rect 55033 -23 55079 23
rect 55157 -23 55203 23
rect 55281 -23 55327 23
rect 55405 -23 55451 23
rect 55529 -23 55575 23
rect 55653 -23 55699 23
rect 55777 -23 55823 23
rect 55901 -23 55947 23
rect 56025 -23 56071 23
rect 56149 -23 56195 23
rect 56273 -23 56319 23
rect 56397 -23 56443 23
rect 56521 -23 56567 23
rect 56645 -23 56691 23
rect 56769 -23 56815 23
rect 56893 -23 56939 23
rect 57017 -23 57063 23
rect 57141 -23 57187 23
rect 57265 -23 57311 23
rect 57389 -23 57435 23
rect 57513 -23 57559 23
rect 57637 -23 57683 23
rect 57761 -23 57807 23
rect 57885 -23 57931 23
rect 58009 -23 58055 23
rect 58133 -23 58179 23
rect 58257 -23 58303 23
rect 58381 -23 58427 23
rect 58505 -23 58551 23
rect 58629 -23 58675 23
rect 58753 -23 58799 23
rect 58877 -23 58923 23
rect 59001 -23 59047 23
rect 59125 -23 59171 23
rect 59249 -23 59295 23
rect 59373 -23 59419 23
rect 59497 -23 59543 23
rect 59621 -23 59667 23
rect 59745 -23 59791 23
rect 59869 -23 59915 23
rect 59993 -23 60039 23
rect 60117 -23 60163 23
rect 60241 -23 60287 23
rect 60365 -23 60411 23
rect 60489 -23 60535 23
rect 60613 -23 60659 23
rect 60737 -23 60783 23
rect 60861 -23 60907 23
rect 60985 -23 61031 23
rect 61109 -23 61155 23
rect 61233 -23 61279 23
rect 61357 -23 61403 23
rect 61481 -23 61527 23
rect 61605 -23 61651 23
rect 61729 -23 61775 23
rect 61853 -23 61899 23
rect 61977 -23 62023 23
rect 62101 -23 62147 23
rect 62225 -23 62271 23
rect 62349 -23 62395 23
rect 62473 -23 62519 23
rect 62597 -23 62643 23
rect 62721 -23 62767 23
rect 62845 -23 62891 23
rect 62969 -23 63015 23
rect 63093 -23 63139 23
rect 63217 -23 63263 23
rect 63341 -23 63387 23
rect 63465 -23 63511 23
rect 63589 -23 63635 23
rect 63713 -23 63759 23
rect 63837 -23 63883 23
rect 63961 -23 64007 23
rect 64085 -23 64131 23
rect 64209 -23 64255 23
rect 64333 -23 64379 23
rect 64457 -23 64503 23
rect 64581 -23 64627 23
rect 64705 -23 64751 23
rect 64829 -23 64875 23
rect 64953 -23 64999 23
rect 65077 -23 65123 23
rect 65201 -23 65247 23
rect 65325 -23 65371 23
rect 65449 -23 65495 23
rect 65573 -23 65619 23
rect 65697 -23 65743 23
rect 65821 -23 65867 23
rect 65945 -23 65991 23
rect 66069 -23 66115 23
rect 66193 -23 66239 23
rect 66317 -23 66363 23
rect 66441 -23 66487 23
rect 66565 -23 66611 23
rect 66689 -23 66735 23
rect 66813 -23 66859 23
rect 66937 -23 66983 23
rect 67061 -23 67107 23
rect 67185 -23 67231 23
rect 67309 -23 67355 23
rect 67433 -23 67479 23
rect 67557 -23 67603 23
rect 67681 -23 67727 23
rect 67805 -23 67851 23
rect 67929 -23 67975 23
rect 68053 -23 68099 23
rect 68177 -23 68223 23
rect 68301 -23 68347 23
rect 68425 -23 68471 23
rect 68549 -23 68595 23
rect 68673 -23 68719 23
rect 68797 -23 68843 23
rect 68921 -23 68967 23
rect 69045 -23 69091 23
rect 69169 -23 69215 23
rect 69293 -23 69339 23
rect 69417 -23 69463 23
rect 69541 -23 69587 23
rect 69665 -23 69711 23
rect 69789 -23 69835 23
rect 69913 -23 69959 23
rect 70037 -23 70083 23
rect 70161 -23 70207 23
rect 70285 -23 70331 23
rect 70409 -23 70455 23
rect 70533 -23 70579 23
rect 70657 -23 70703 23
rect 70781 -23 70827 23
rect 70905 -23 70951 23
rect 71029 -23 71075 23
rect 71153 -23 71199 23
rect 71277 -23 71323 23
rect 71401 -23 71447 23
rect 71525 -23 71571 23
rect 71649 -23 71695 23
rect 71773 -23 71819 23
rect 71897 -23 71943 23
rect 72021 -23 72067 23
rect 72145 -23 72191 23
rect 72269 -23 72315 23
rect 72393 -23 72439 23
rect 72517 -23 72563 23
rect 72641 -23 72687 23
rect 72765 -23 72811 23
rect 72889 -23 72935 23
rect 73013 -23 73059 23
rect 73137 -23 73183 23
rect 73261 -23 73307 23
rect 73385 -23 73431 23
rect 73509 -23 73555 23
rect 73633 -23 73679 23
rect 73757 -23 73803 23
rect 73881 -23 73927 23
rect 74005 -23 74051 23
rect 74129 -23 74175 23
rect 74253 -23 74299 23
rect 74377 -23 74423 23
rect 74501 -23 74547 23
rect 74625 -23 74671 23
rect 74749 -23 74795 23
rect 74873 -23 74919 23
rect 74997 -23 75043 23
rect 75121 -23 75167 23
rect 75245 -23 75291 23
rect 75369 -23 75415 23
rect 75493 -23 75539 23
rect 75617 -23 75663 23
rect 75741 -23 75787 23
rect 75865 -23 75911 23
rect 75989 -23 76035 23
rect 76113 -23 76159 23
rect 76237 -23 76283 23
rect 76361 -23 76407 23
rect 76485 -23 76531 23
rect 76609 -23 76655 23
rect 76733 -23 76779 23
rect 76857 -23 76903 23
rect 76981 -23 77027 23
rect 77105 -23 77151 23
rect 77229 -23 77275 23
rect 77353 -23 77399 23
rect 77477 -23 77523 23
rect 77601 -23 77647 23
rect 77725 -23 77771 23
rect 77849 -23 77895 23
rect 77973 -23 78019 23
rect 78097 -23 78143 23
rect 78221 -23 78267 23
rect 78345 -23 78391 23
rect 78469 -23 78515 23
rect 78593 -23 78639 23
rect 78717 -23 78763 23
rect 78841 -23 78887 23
rect 78965 -23 79011 23
rect 79089 -23 79135 23
rect 79213 -23 79259 23
rect 79337 -23 79383 23
rect 79461 -23 79507 23
rect 79585 -23 79631 23
rect 79709 -23 79755 23
rect 79833 -23 79879 23
rect 79957 -23 80003 23
rect 80081 -23 80127 23
rect 80205 -23 80251 23
rect 80329 -23 80375 23
rect 80453 -23 80499 23
rect 80577 -23 80623 23
rect 80701 -23 80747 23
rect 80825 -23 80871 23
rect 80949 -23 80995 23
rect 81073 -23 81119 23
rect 81197 -23 81243 23
rect 81321 -23 81367 23
rect 81445 -23 81491 23
rect 81569 -23 81615 23
rect 81693 -23 81739 23
rect 81817 -23 81863 23
rect 81941 -23 81987 23
rect 82065 -23 82111 23
rect 82189 -23 82235 23
rect 82313 -23 82359 23
rect 82437 -23 82483 23
rect 82561 -23 82607 23
rect 82685 -23 82731 23
rect 82809 -23 82855 23
rect 82933 -23 82979 23
rect 83057 -23 83103 23
rect 83181 -23 83227 23
rect 83305 -23 83351 23
rect 83429 -23 83475 23
rect 83553 -23 83599 23
rect 83677 -23 83723 23
rect 83801 -23 83847 23
rect 83925 -23 83971 23
rect 84049 -23 84095 23
rect 84173 -23 84219 23
rect 84297 -23 84343 23
rect 84421 -23 84467 23
rect 84545 -23 84591 23
rect 84669 -23 84715 23
rect 84793 -23 84839 23
rect 84917 -23 84963 23
rect 85041 -23 85087 23
rect 85165 -23 85211 23
rect 85289 -23 85335 23
rect 85413 -23 85459 23
rect 85537 -23 85583 23
<< metal1 >>
rect -34 395 85594 406
rect -34 349 -23 395
rect 23 349 101 395
rect 147 349 225 395
rect 271 349 349 395
rect 395 349 473 395
rect 519 349 597 395
rect 643 349 721 395
rect 767 349 845 395
rect 891 349 969 395
rect 1015 349 1093 395
rect 1139 349 1217 395
rect 1263 349 1341 395
rect 1387 349 1465 395
rect 1511 349 1589 395
rect 1635 349 1713 395
rect 1759 349 1837 395
rect 1883 349 1961 395
rect 2007 349 2085 395
rect 2131 349 2209 395
rect 2255 349 2333 395
rect 2379 349 2457 395
rect 2503 349 2581 395
rect 2627 349 2705 395
rect 2751 349 2829 395
rect 2875 349 2953 395
rect 2999 349 3077 395
rect 3123 349 3201 395
rect 3247 349 3325 395
rect 3371 349 3449 395
rect 3495 349 3573 395
rect 3619 349 3697 395
rect 3743 349 3821 395
rect 3867 349 3945 395
rect 3991 349 4069 395
rect 4115 349 4193 395
rect 4239 349 4317 395
rect 4363 349 4441 395
rect 4487 349 4565 395
rect 4611 349 4689 395
rect 4735 349 4813 395
rect 4859 349 4937 395
rect 4983 349 5061 395
rect 5107 349 5185 395
rect 5231 349 5309 395
rect 5355 349 5433 395
rect 5479 349 5557 395
rect 5603 349 5681 395
rect 5727 349 5805 395
rect 5851 349 5929 395
rect 5975 349 6053 395
rect 6099 349 6177 395
rect 6223 349 6301 395
rect 6347 349 6425 395
rect 6471 349 6549 395
rect 6595 349 6673 395
rect 6719 349 6797 395
rect 6843 349 6921 395
rect 6967 349 7045 395
rect 7091 349 7169 395
rect 7215 349 7293 395
rect 7339 349 7417 395
rect 7463 349 7541 395
rect 7587 349 7665 395
rect 7711 349 7789 395
rect 7835 349 7913 395
rect 7959 349 8037 395
rect 8083 349 8161 395
rect 8207 349 8285 395
rect 8331 349 8409 395
rect 8455 349 8533 395
rect 8579 349 8657 395
rect 8703 349 8781 395
rect 8827 349 8905 395
rect 8951 349 9029 395
rect 9075 349 9153 395
rect 9199 349 9277 395
rect 9323 349 9401 395
rect 9447 349 9525 395
rect 9571 349 9649 395
rect 9695 349 9773 395
rect 9819 349 9897 395
rect 9943 349 10021 395
rect 10067 349 10145 395
rect 10191 349 10269 395
rect 10315 349 10393 395
rect 10439 349 10517 395
rect 10563 349 10641 395
rect 10687 349 10765 395
rect 10811 349 10889 395
rect 10935 349 11013 395
rect 11059 349 11137 395
rect 11183 349 11261 395
rect 11307 349 11385 395
rect 11431 349 11509 395
rect 11555 349 11633 395
rect 11679 349 11757 395
rect 11803 349 11881 395
rect 11927 349 12005 395
rect 12051 349 12129 395
rect 12175 349 12253 395
rect 12299 349 12377 395
rect 12423 349 12501 395
rect 12547 349 12625 395
rect 12671 349 12749 395
rect 12795 349 12873 395
rect 12919 349 12997 395
rect 13043 349 13121 395
rect 13167 349 13245 395
rect 13291 349 13369 395
rect 13415 349 13493 395
rect 13539 349 13617 395
rect 13663 349 13741 395
rect 13787 349 13865 395
rect 13911 349 13989 395
rect 14035 349 14113 395
rect 14159 349 14237 395
rect 14283 349 14361 395
rect 14407 349 14485 395
rect 14531 349 14609 395
rect 14655 349 14733 395
rect 14779 349 14857 395
rect 14903 349 14981 395
rect 15027 349 15105 395
rect 15151 349 15229 395
rect 15275 349 15353 395
rect 15399 349 15477 395
rect 15523 349 15601 395
rect 15647 349 15725 395
rect 15771 349 15849 395
rect 15895 349 15973 395
rect 16019 349 16097 395
rect 16143 349 16221 395
rect 16267 349 16345 395
rect 16391 349 16469 395
rect 16515 349 16593 395
rect 16639 349 16717 395
rect 16763 349 16841 395
rect 16887 349 16965 395
rect 17011 349 17089 395
rect 17135 349 17213 395
rect 17259 349 17337 395
rect 17383 349 17461 395
rect 17507 349 17585 395
rect 17631 349 17709 395
rect 17755 349 17833 395
rect 17879 349 17957 395
rect 18003 349 18081 395
rect 18127 349 18205 395
rect 18251 349 18329 395
rect 18375 349 18453 395
rect 18499 349 18577 395
rect 18623 349 18701 395
rect 18747 349 18825 395
rect 18871 349 18949 395
rect 18995 349 19073 395
rect 19119 349 19197 395
rect 19243 349 19321 395
rect 19367 349 19445 395
rect 19491 349 19569 395
rect 19615 349 19693 395
rect 19739 349 19817 395
rect 19863 349 19941 395
rect 19987 349 20065 395
rect 20111 349 20189 395
rect 20235 349 20313 395
rect 20359 349 20437 395
rect 20483 349 20561 395
rect 20607 349 20685 395
rect 20731 349 20809 395
rect 20855 349 20933 395
rect 20979 349 21057 395
rect 21103 349 21181 395
rect 21227 349 21305 395
rect 21351 349 21429 395
rect 21475 349 21553 395
rect 21599 349 21677 395
rect 21723 349 21801 395
rect 21847 349 21925 395
rect 21971 349 22049 395
rect 22095 349 22173 395
rect 22219 349 22297 395
rect 22343 349 22421 395
rect 22467 349 22545 395
rect 22591 349 22669 395
rect 22715 349 22793 395
rect 22839 349 22917 395
rect 22963 349 23041 395
rect 23087 349 23165 395
rect 23211 349 23289 395
rect 23335 349 23413 395
rect 23459 349 23537 395
rect 23583 349 23661 395
rect 23707 349 23785 395
rect 23831 349 23909 395
rect 23955 349 24033 395
rect 24079 349 24157 395
rect 24203 349 24281 395
rect 24327 349 24405 395
rect 24451 349 24529 395
rect 24575 349 24653 395
rect 24699 349 24777 395
rect 24823 349 24901 395
rect 24947 349 25025 395
rect 25071 349 25149 395
rect 25195 349 25273 395
rect 25319 349 25397 395
rect 25443 349 25521 395
rect 25567 349 25645 395
rect 25691 349 25769 395
rect 25815 349 25893 395
rect 25939 349 26017 395
rect 26063 349 26141 395
rect 26187 349 26265 395
rect 26311 349 26389 395
rect 26435 349 26513 395
rect 26559 349 26637 395
rect 26683 349 26761 395
rect 26807 349 26885 395
rect 26931 349 27009 395
rect 27055 349 27133 395
rect 27179 349 27257 395
rect 27303 349 27381 395
rect 27427 349 27505 395
rect 27551 349 27629 395
rect 27675 349 27753 395
rect 27799 349 27877 395
rect 27923 349 28001 395
rect 28047 349 28125 395
rect 28171 349 28249 395
rect 28295 349 28373 395
rect 28419 349 28497 395
rect 28543 349 28621 395
rect 28667 349 28745 395
rect 28791 349 28869 395
rect 28915 349 28993 395
rect 29039 349 29117 395
rect 29163 349 29241 395
rect 29287 349 29365 395
rect 29411 349 29489 395
rect 29535 349 29613 395
rect 29659 349 29737 395
rect 29783 349 29861 395
rect 29907 349 29985 395
rect 30031 349 30109 395
rect 30155 349 30233 395
rect 30279 349 30357 395
rect 30403 349 30481 395
rect 30527 349 30605 395
rect 30651 349 30729 395
rect 30775 349 30853 395
rect 30899 349 30977 395
rect 31023 349 31101 395
rect 31147 349 31225 395
rect 31271 349 31349 395
rect 31395 349 31473 395
rect 31519 349 31597 395
rect 31643 349 31721 395
rect 31767 349 31845 395
rect 31891 349 31969 395
rect 32015 349 32093 395
rect 32139 349 32217 395
rect 32263 349 32341 395
rect 32387 349 32465 395
rect 32511 349 32589 395
rect 32635 349 32713 395
rect 32759 349 32837 395
rect 32883 349 32961 395
rect 33007 349 33085 395
rect 33131 349 33209 395
rect 33255 349 33333 395
rect 33379 349 33457 395
rect 33503 349 33581 395
rect 33627 349 33705 395
rect 33751 349 33829 395
rect 33875 349 33953 395
rect 33999 349 34077 395
rect 34123 349 34201 395
rect 34247 349 34325 395
rect 34371 349 34449 395
rect 34495 349 34573 395
rect 34619 349 34697 395
rect 34743 349 34821 395
rect 34867 349 34945 395
rect 34991 349 35069 395
rect 35115 349 35193 395
rect 35239 349 35317 395
rect 35363 349 35441 395
rect 35487 349 35565 395
rect 35611 349 35689 395
rect 35735 349 35813 395
rect 35859 349 35937 395
rect 35983 349 36061 395
rect 36107 349 36185 395
rect 36231 349 36309 395
rect 36355 349 36433 395
rect 36479 349 36557 395
rect 36603 349 36681 395
rect 36727 349 36805 395
rect 36851 349 36929 395
rect 36975 349 37053 395
rect 37099 349 37177 395
rect 37223 349 37301 395
rect 37347 349 37425 395
rect 37471 349 37549 395
rect 37595 349 37673 395
rect 37719 349 37797 395
rect 37843 349 37921 395
rect 37967 349 38045 395
rect 38091 349 38169 395
rect 38215 349 38293 395
rect 38339 349 38417 395
rect 38463 349 38541 395
rect 38587 349 38665 395
rect 38711 349 38789 395
rect 38835 349 38913 395
rect 38959 349 39037 395
rect 39083 349 39161 395
rect 39207 349 39285 395
rect 39331 349 39409 395
rect 39455 349 39533 395
rect 39579 349 39657 395
rect 39703 349 39781 395
rect 39827 349 39905 395
rect 39951 349 40029 395
rect 40075 349 40153 395
rect 40199 349 40277 395
rect 40323 349 40401 395
rect 40447 349 40525 395
rect 40571 349 40649 395
rect 40695 349 40773 395
rect 40819 349 40897 395
rect 40943 349 41021 395
rect 41067 349 41145 395
rect 41191 349 41269 395
rect 41315 349 41393 395
rect 41439 349 41517 395
rect 41563 349 41641 395
rect 41687 349 41765 395
rect 41811 349 41889 395
rect 41935 349 42013 395
rect 42059 349 42137 395
rect 42183 349 42261 395
rect 42307 349 42385 395
rect 42431 349 42509 395
rect 42555 349 42633 395
rect 42679 349 42757 395
rect 42803 349 42881 395
rect 42927 349 43005 395
rect 43051 349 43129 395
rect 43175 349 43253 395
rect 43299 349 43377 395
rect 43423 349 43501 395
rect 43547 349 43625 395
rect 43671 349 43749 395
rect 43795 349 43873 395
rect 43919 349 43997 395
rect 44043 349 44121 395
rect 44167 349 44245 395
rect 44291 349 44369 395
rect 44415 349 44493 395
rect 44539 349 44617 395
rect 44663 349 44741 395
rect 44787 349 44865 395
rect 44911 349 44989 395
rect 45035 349 45113 395
rect 45159 349 45237 395
rect 45283 349 45361 395
rect 45407 349 45485 395
rect 45531 349 45609 395
rect 45655 349 45733 395
rect 45779 349 45857 395
rect 45903 349 45981 395
rect 46027 349 46105 395
rect 46151 349 46229 395
rect 46275 349 46353 395
rect 46399 349 46477 395
rect 46523 349 46601 395
rect 46647 349 46725 395
rect 46771 349 46849 395
rect 46895 349 46973 395
rect 47019 349 47097 395
rect 47143 349 47221 395
rect 47267 349 47345 395
rect 47391 349 47469 395
rect 47515 349 47593 395
rect 47639 349 47717 395
rect 47763 349 47841 395
rect 47887 349 47965 395
rect 48011 349 48089 395
rect 48135 349 48213 395
rect 48259 349 48337 395
rect 48383 349 48461 395
rect 48507 349 48585 395
rect 48631 349 48709 395
rect 48755 349 48833 395
rect 48879 349 48957 395
rect 49003 349 49081 395
rect 49127 349 49205 395
rect 49251 349 49329 395
rect 49375 349 49453 395
rect 49499 349 49577 395
rect 49623 349 49701 395
rect 49747 349 49825 395
rect 49871 349 49949 395
rect 49995 349 50073 395
rect 50119 349 50197 395
rect 50243 349 50321 395
rect 50367 349 50445 395
rect 50491 349 50569 395
rect 50615 349 50693 395
rect 50739 349 50817 395
rect 50863 349 50941 395
rect 50987 349 51065 395
rect 51111 349 51189 395
rect 51235 349 51313 395
rect 51359 349 51437 395
rect 51483 349 51561 395
rect 51607 349 51685 395
rect 51731 349 51809 395
rect 51855 349 51933 395
rect 51979 349 52057 395
rect 52103 349 52181 395
rect 52227 349 52305 395
rect 52351 349 52429 395
rect 52475 349 52553 395
rect 52599 349 52677 395
rect 52723 349 52801 395
rect 52847 349 52925 395
rect 52971 349 53049 395
rect 53095 349 53173 395
rect 53219 349 53297 395
rect 53343 349 53421 395
rect 53467 349 53545 395
rect 53591 349 53669 395
rect 53715 349 53793 395
rect 53839 349 53917 395
rect 53963 349 54041 395
rect 54087 349 54165 395
rect 54211 349 54289 395
rect 54335 349 54413 395
rect 54459 349 54537 395
rect 54583 349 54661 395
rect 54707 349 54785 395
rect 54831 349 54909 395
rect 54955 349 55033 395
rect 55079 349 55157 395
rect 55203 349 55281 395
rect 55327 349 55405 395
rect 55451 349 55529 395
rect 55575 349 55653 395
rect 55699 349 55777 395
rect 55823 349 55901 395
rect 55947 349 56025 395
rect 56071 349 56149 395
rect 56195 349 56273 395
rect 56319 349 56397 395
rect 56443 349 56521 395
rect 56567 349 56645 395
rect 56691 349 56769 395
rect 56815 349 56893 395
rect 56939 349 57017 395
rect 57063 349 57141 395
rect 57187 349 57265 395
rect 57311 349 57389 395
rect 57435 349 57513 395
rect 57559 349 57637 395
rect 57683 349 57761 395
rect 57807 349 57885 395
rect 57931 349 58009 395
rect 58055 349 58133 395
rect 58179 349 58257 395
rect 58303 349 58381 395
rect 58427 349 58505 395
rect 58551 349 58629 395
rect 58675 349 58753 395
rect 58799 349 58877 395
rect 58923 349 59001 395
rect 59047 349 59125 395
rect 59171 349 59249 395
rect 59295 349 59373 395
rect 59419 349 59497 395
rect 59543 349 59621 395
rect 59667 349 59745 395
rect 59791 349 59869 395
rect 59915 349 59993 395
rect 60039 349 60117 395
rect 60163 349 60241 395
rect 60287 349 60365 395
rect 60411 349 60489 395
rect 60535 349 60613 395
rect 60659 349 60737 395
rect 60783 349 60861 395
rect 60907 349 60985 395
rect 61031 349 61109 395
rect 61155 349 61233 395
rect 61279 349 61357 395
rect 61403 349 61481 395
rect 61527 349 61605 395
rect 61651 349 61729 395
rect 61775 349 61853 395
rect 61899 349 61977 395
rect 62023 349 62101 395
rect 62147 349 62225 395
rect 62271 349 62349 395
rect 62395 349 62473 395
rect 62519 349 62597 395
rect 62643 349 62721 395
rect 62767 349 62845 395
rect 62891 349 62969 395
rect 63015 349 63093 395
rect 63139 349 63217 395
rect 63263 349 63341 395
rect 63387 349 63465 395
rect 63511 349 63589 395
rect 63635 349 63713 395
rect 63759 349 63837 395
rect 63883 349 63961 395
rect 64007 349 64085 395
rect 64131 349 64209 395
rect 64255 349 64333 395
rect 64379 349 64457 395
rect 64503 349 64581 395
rect 64627 349 64705 395
rect 64751 349 64829 395
rect 64875 349 64953 395
rect 64999 349 65077 395
rect 65123 349 65201 395
rect 65247 349 65325 395
rect 65371 349 65449 395
rect 65495 349 65573 395
rect 65619 349 65697 395
rect 65743 349 65821 395
rect 65867 349 65945 395
rect 65991 349 66069 395
rect 66115 349 66193 395
rect 66239 349 66317 395
rect 66363 349 66441 395
rect 66487 349 66565 395
rect 66611 349 66689 395
rect 66735 349 66813 395
rect 66859 349 66937 395
rect 66983 349 67061 395
rect 67107 349 67185 395
rect 67231 349 67309 395
rect 67355 349 67433 395
rect 67479 349 67557 395
rect 67603 349 67681 395
rect 67727 349 67805 395
rect 67851 349 67929 395
rect 67975 349 68053 395
rect 68099 349 68177 395
rect 68223 349 68301 395
rect 68347 349 68425 395
rect 68471 349 68549 395
rect 68595 349 68673 395
rect 68719 349 68797 395
rect 68843 349 68921 395
rect 68967 349 69045 395
rect 69091 349 69169 395
rect 69215 349 69293 395
rect 69339 349 69417 395
rect 69463 349 69541 395
rect 69587 349 69665 395
rect 69711 349 69789 395
rect 69835 349 69913 395
rect 69959 349 70037 395
rect 70083 349 70161 395
rect 70207 349 70285 395
rect 70331 349 70409 395
rect 70455 349 70533 395
rect 70579 349 70657 395
rect 70703 349 70781 395
rect 70827 349 70905 395
rect 70951 349 71029 395
rect 71075 349 71153 395
rect 71199 349 71277 395
rect 71323 349 71401 395
rect 71447 349 71525 395
rect 71571 349 71649 395
rect 71695 349 71773 395
rect 71819 349 71897 395
rect 71943 349 72021 395
rect 72067 349 72145 395
rect 72191 349 72269 395
rect 72315 349 72393 395
rect 72439 349 72517 395
rect 72563 349 72641 395
rect 72687 349 72765 395
rect 72811 349 72889 395
rect 72935 349 73013 395
rect 73059 349 73137 395
rect 73183 349 73261 395
rect 73307 349 73385 395
rect 73431 349 73509 395
rect 73555 349 73633 395
rect 73679 349 73757 395
rect 73803 349 73881 395
rect 73927 349 74005 395
rect 74051 349 74129 395
rect 74175 349 74253 395
rect 74299 349 74377 395
rect 74423 349 74501 395
rect 74547 349 74625 395
rect 74671 349 74749 395
rect 74795 349 74873 395
rect 74919 349 74997 395
rect 75043 349 75121 395
rect 75167 349 75245 395
rect 75291 349 75369 395
rect 75415 349 75493 395
rect 75539 349 75617 395
rect 75663 349 75741 395
rect 75787 349 75865 395
rect 75911 349 75989 395
rect 76035 349 76113 395
rect 76159 349 76237 395
rect 76283 349 76361 395
rect 76407 349 76485 395
rect 76531 349 76609 395
rect 76655 349 76733 395
rect 76779 349 76857 395
rect 76903 349 76981 395
rect 77027 349 77105 395
rect 77151 349 77229 395
rect 77275 349 77353 395
rect 77399 349 77477 395
rect 77523 349 77601 395
rect 77647 349 77725 395
rect 77771 349 77849 395
rect 77895 349 77973 395
rect 78019 349 78097 395
rect 78143 349 78221 395
rect 78267 349 78345 395
rect 78391 349 78469 395
rect 78515 349 78593 395
rect 78639 349 78717 395
rect 78763 349 78841 395
rect 78887 349 78965 395
rect 79011 349 79089 395
rect 79135 349 79213 395
rect 79259 349 79337 395
rect 79383 349 79461 395
rect 79507 349 79585 395
rect 79631 349 79709 395
rect 79755 349 79833 395
rect 79879 349 79957 395
rect 80003 349 80081 395
rect 80127 349 80205 395
rect 80251 349 80329 395
rect 80375 349 80453 395
rect 80499 349 80577 395
rect 80623 349 80701 395
rect 80747 349 80825 395
rect 80871 349 80949 395
rect 80995 349 81073 395
rect 81119 349 81197 395
rect 81243 349 81321 395
rect 81367 349 81445 395
rect 81491 349 81569 395
rect 81615 349 81693 395
rect 81739 349 81817 395
rect 81863 349 81941 395
rect 81987 349 82065 395
rect 82111 349 82189 395
rect 82235 349 82313 395
rect 82359 349 82437 395
rect 82483 349 82561 395
rect 82607 349 82685 395
rect 82731 349 82809 395
rect 82855 349 82933 395
rect 82979 349 83057 395
rect 83103 349 83181 395
rect 83227 349 83305 395
rect 83351 349 83429 395
rect 83475 349 83553 395
rect 83599 349 83677 395
rect 83723 349 83801 395
rect 83847 349 83925 395
rect 83971 349 84049 395
rect 84095 349 84173 395
rect 84219 349 84297 395
rect 84343 349 84421 395
rect 84467 349 84545 395
rect 84591 349 84669 395
rect 84715 349 84793 395
rect 84839 349 84917 395
rect 84963 349 85041 395
rect 85087 349 85165 395
rect 85211 349 85289 395
rect 85335 349 85413 395
rect 85459 349 85537 395
rect 85583 349 85594 395
rect -34 271 85594 349
rect -34 225 -23 271
rect 23 225 101 271
rect 147 225 225 271
rect 271 225 349 271
rect 395 225 473 271
rect 519 225 597 271
rect 643 225 721 271
rect 767 225 845 271
rect 891 225 969 271
rect 1015 225 1093 271
rect 1139 225 1217 271
rect 1263 225 1341 271
rect 1387 225 1465 271
rect 1511 225 1589 271
rect 1635 225 1713 271
rect 1759 225 1837 271
rect 1883 225 1961 271
rect 2007 225 2085 271
rect 2131 225 2209 271
rect 2255 225 2333 271
rect 2379 225 2457 271
rect 2503 225 2581 271
rect 2627 225 2705 271
rect 2751 225 2829 271
rect 2875 225 2953 271
rect 2999 225 3077 271
rect 3123 225 3201 271
rect 3247 225 3325 271
rect 3371 225 3449 271
rect 3495 225 3573 271
rect 3619 225 3697 271
rect 3743 225 3821 271
rect 3867 225 3945 271
rect 3991 225 4069 271
rect 4115 225 4193 271
rect 4239 225 4317 271
rect 4363 225 4441 271
rect 4487 225 4565 271
rect 4611 225 4689 271
rect 4735 225 4813 271
rect 4859 225 4937 271
rect 4983 225 5061 271
rect 5107 225 5185 271
rect 5231 225 5309 271
rect 5355 225 5433 271
rect 5479 225 5557 271
rect 5603 225 5681 271
rect 5727 225 5805 271
rect 5851 225 5929 271
rect 5975 225 6053 271
rect 6099 225 6177 271
rect 6223 225 6301 271
rect 6347 225 6425 271
rect 6471 225 6549 271
rect 6595 225 6673 271
rect 6719 225 6797 271
rect 6843 225 6921 271
rect 6967 225 7045 271
rect 7091 225 7169 271
rect 7215 225 7293 271
rect 7339 225 7417 271
rect 7463 225 7541 271
rect 7587 225 7665 271
rect 7711 225 7789 271
rect 7835 225 7913 271
rect 7959 225 8037 271
rect 8083 225 8161 271
rect 8207 225 8285 271
rect 8331 225 8409 271
rect 8455 225 8533 271
rect 8579 225 8657 271
rect 8703 225 8781 271
rect 8827 225 8905 271
rect 8951 225 9029 271
rect 9075 225 9153 271
rect 9199 225 9277 271
rect 9323 225 9401 271
rect 9447 225 9525 271
rect 9571 225 9649 271
rect 9695 225 9773 271
rect 9819 225 9897 271
rect 9943 225 10021 271
rect 10067 225 10145 271
rect 10191 225 10269 271
rect 10315 225 10393 271
rect 10439 225 10517 271
rect 10563 225 10641 271
rect 10687 225 10765 271
rect 10811 225 10889 271
rect 10935 225 11013 271
rect 11059 225 11137 271
rect 11183 225 11261 271
rect 11307 225 11385 271
rect 11431 225 11509 271
rect 11555 225 11633 271
rect 11679 225 11757 271
rect 11803 225 11881 271
rect 11927 225 12005 271
rect 12051 225 12129 271
rect 12175 225 12253 271
rect 12299 225 12377 271
rect 12423 225 12501 271
rect 12547 225 12625 271
rect 12671 225 12749 271
rect 12795 225 12873 271
rect 12919 225 12997 271
rect 13043 225 13121 271
rect 13167 225 13245 271
rect 13291 225 13369 271
rect 13415 225 13493 271
rect 13539 225 13617 271
rect 13663 225 13741 271
rect 13787 225 13865 271
rect 13911 225 13989 271
rect 14035 225 14113 271
rect 14159 225 14237 271
rect 14283 225 14361 271
rect 14407 225 14485 271
rect 14531 225 14609 271
rect 14655 225 14733 271
rect 14779 225 14857 271
rect 14903 225 14981 271
rect 15027 225 15105 271
rect 15151 225 15229 271
rect 15275 225 15353 271
rect 15399 225 15477 271
rect 15523 225 15601 271
rect 15647 225 15725 271
rect 15771 225 15849 271
rect 15895 225 15973 271
rect 16019 225 16097 271
rect 16143 225 16221 271
rect 16267 225 16345 271
rect 16391 225 16469 271
rect 16515 225 16593 271
rect 16639 225 16717 271
rect 16763 225 16841 271
rect 16887 225 16965 271
rect 17011 225 17089 271
rect 17135 225 17213 271
rect 17259 225 17337 271
rect 17383 225 17461 271
rect 17507 225 17585 271
rect 17631 225 17709 271
rect 17755 225 17833 271
rect 17879 225 17957 271
rect 18003 225 18081 271
rect 18127 225 18205 271
rect 18251 225 18329 271
rect 18375 225 18453 271
rect 18499 225 18577 271
rect 18623 225 18701 271
rect 18747 225 18825 271
rect 18871 225 18949 271
rect 18995 225 19073 271
rect 19119 225 19197 271
rect 19243 225 19321 271
rect 19367 225 19445 271
rect 19491 225 19569 271
rect 19615 225 19693 271
rect 19739 225 19817 271
rect 19863 225 19941 271
rect 19987 225 20065 271
rect 20111 225 20189 271
rect 20235 225 20313 271
rect 20359 225 20437 271
rect 20483 225 20561 271
rect 20607 225 20685 271
rect 20731 225 20809 271
rect 20855 225 20933 271
rect 20979 225 21057 271
rect 21103 225 21181 271
rect 21227 225 21305 271
rect 21351 225 21429 271
rect 21475 225 21553 271
rect 21599 225 21677 271
rect 21723 225 21801 271
rect 21847 225 21925 271
rect 21971 225 22049 271
rect 22095 225 22173 271
rect 22219 225 22297 271
rect 22343 225 22421 271
rect 22467 225 22545 271
rect 22591 225 22669 271
rect 22715 225 22793 271
rect 22839 225 22917 271
rect 22963 225 23041 271
rect 23087 225 23165 271
rect 23211 225 23289 271
rect 23335 225 23413 271
rect 23459 225 23537 271
rect 23583 225 23661 271
rect 23707 225 23785 271
rect 23831 225 23909 271
rect 23955 225 24033 271
rect 24079 225 24157 271
rect 24203 225 24281 271
rect 24327 225 24405 271
rect 24451 225 24529 271
rect 24575 225 24653 271
rect 24699 225 24777 271
rect 24823 225 24901 271
rect 24947 225 25025 271
rect 25071 225 25149 271
rect 25195 225 25273 271
rect 25319 225 25397 271
rect 25443 225 25521 271
rect 25567 225 25645 271
rect 25691 225 25769 271
rect 25815 225 25893 271
rect 25939 225 26017 271
rect 26063 225 26141 271
rect 26187 225 26265 271
rect 26311 225 26389 271
rect 26435 225 26513 271
rect 26559 225 26637 271
rect 26683 225 26761 271
rect 26807 225 26885 271
rect 26931 225 27009 271
rect 27055 225 27133 271
rect 27179 225 27257 271
rect 27303 225 27381 271
rect 27427 225 27505 271
rect 27551 225 27629 271
rect 27675 225 27753 271
rect 27799 225 27877 271
rect 27923 225 28001 271
rect 28047 225 28125 271
rect 28171 225 28249 271
rect 28295 225 28373 271
rect 28419 225 28497 271
rect 28543 225 28621 271
rect 28667 225 28745 271
rect 28791 225 28869 271
rect 28915 225 28993 271
rect 29039 225 29117 271
rect 29163 225 29241 271
rect 29287 225 29365 271
rect 29411 225 29489 271
rect 29535 225 29613 271
rect 29659 225 29737 271
rect 29783 225 29861 271
rect 29907 225 29985 271
rect 30031 225 30109 271
rect 30155 225 30233 271
rect 30279 225 30357 271
rect 30403 225 30481 271
rect 30527 225 30605 271
rect 30651 225 30729 271
rect 30775 225 30853 271
rect 30899 225 30977 271
rect 31023 225 31101 271
rect 31147 225 31225 271
rect 31271 225 31349 271
rect 31395 225 31473 271
rect 31519 225 31597 271
rect 31643 225 31721 271
rect 31767 225 31845 271
rect 31891 225 31969 271
rect 32015 225 32093 271
rect 32139 225 32217 271
rect 32263 225 32341 271
rect 32387 225 32465 271
rect 32511 225 32589 271
rect 32635 225 32713 271
rect 32759 225 32837 271
rect 32883 225 32961 271
rect 33007 225 33085 271
rect 33131 225 33209 271
rect 33255 225 33333 271
rect 33379 225 33457 271
rect 33503 225 33581 271
rect 33627 225 33705 271
rect 33751 225 33829 271
rect 33875 225 33953 271
rect 33999 225 34077 271
rect 34123 225 34201 271
rect 34247 225 34325 271
rect 34371 225 34449 271
rect 34495 225 34573 271
rect 34619 225 34697 271
rect 34743 225 34821 271
rect 34867 225 34945 271
rect 34991 225 35069 271
rect 35115 225 35193 271
rect 35239 225 35317 271
rect 35363 225 35441 271
rect 35487 225 35565 271
rect 35611 225 35689 271
rect 35735 225 35813 271
rect 35859 225 35937 271
rect 35983 225 36061 271
rect 36107 225 36185 271
rect 36231 225 36309 271
rect 36355 225 36433 271
rect 36479 225 36557 271
rect 36603 225 36681 271
rect 36727 225 36805 271
rect 36851 225 36929 271
rect 36975 225 37053 271
rect 37099 225 37177 271
rect 37223 225 37301 271
rect 37347 225 37425 271
rect 37471 225 37549 271
rect 37595 225 37673 271
rect 37719 225 37797 271
rect 37843 225 37921 271
rect 37967 225 38045 271
rect 38091 225 38169 271
rect 38215 225 38293 271
rect 38339 225 38417 271
rect 38463 225 38541 271
rect 38587 225 38665 271
rect 38711 225 38789 271
rect 38835 225 38913 271
rect 38959 225 39037 271
rect 39083 225 39161 271
rect 39207 225 39285 271
rect 39331 225 39409 271
rect 39455 225 39533 271
rect 39579 225 39657 271
rect 39703 225 39781 271
rect 39827 225 39905 271
rect 39951 225 40029 271
rect 40075 225 40153 271
rect 40199 225 40277 271
rect 40323 225 40401 271
rect 40447 225 40525 271
rect 40571 225 40649 271
rect 40695 225 40773 271
rect 40819 225 40897 271
rect 40943 225 41021 271
rect 41067 225 41145 271
rect 41191 225 41269 271
rect 41315 225 41393 271
rect 41439 225 41517 271
rect 41563 225 41641 271
rect 41687 225 41765 271
rect 41811 225 41889 271
rect 41935 225 42013 271
rect 42059 225 42137 271
rect 42183 225 42261 271
rect 42307 225 42385 271
rect 42431 225 42509 271
rect 42555 225 42633 271
rect 42679 225 42757 271
rect 42803 225 42881 271
rect 42927 225 43005 271
rect 43051 225 43129 271
rect 43175 225 43253 271
rect 43299 225 43377 271
rect 43423 225 43501 271
rect 43547 225 43625 271
rect 43671 225 43749 271
rect 43795 225 43873 271
rect 43919 225 43997 271
rect 44043 225 44121 271
rect 44167 225 44245 271
rect 44291 225 44369 271
rect 44415 225 44493 271
rect 44539 225 44617 271
rect 44663 225 44741 271
rect 44787 225 44865 271
rect 44911 225 44989 271
rect 45035 225 45113 271
rect 45159 225 45237 271
rect 45283 225 45361 271
rect 45407 225 45485 271
rect 45531 225 45609 271
rect 45655 225 45733 271
rect 45779 225 45857 271
rect 45903 225 45981 271
rect 46027 225 46105 271
rect 46151 225 46229 271
rect 46275 225 46353 271
rect 46399 225 46477 271
rect 46523 225 46601 271
rect 46647 225 46725 271
rect 46771 225 46849 271
rect 46895 225 46973 271
rect 47019 225 47097 271
rect 47143 225 47221 271
rect 47267 225 47345 271
rect 47391 225 47469 271
rect 47515 225 47593 271
rect 47639 225 47717 271
rect 47763 225 47841 271
rect 47887 225 47965 271
rect 48011 225 48089 271
rect 48135 225 48213 271
rect 48259 225 48337 271
rect 48383 225 48461 271
rect 48507 225 48585 271
rect 48631 225 48709 271
rect 48755 225 48833 271
rect 48879 225 48957 271
rect 49003 225 49081 271
rect 49127 225 49205 271
rect 49251 225 49329 271
rect 49375 225 49453 271
rect 49499 225 49577 271
rect 49623 225 49701 271
rect 49747 225 49825 271
rect 49871 225 49949 271
rect 49995 225 50073 271
rect 50119 225 50197 271
rect 50243 225 50321 271
rect 50367 225 50445 271
rect 50491 225 50569 271
rect 50615 225 50693 271
rect 50739 225 50817 271
rect 50863 225 50941 271
rect 50987 225 51065 271
rect 51111 225 51189 271
rect 51235 225 51313 271
rect 51359 225 51437 271
rect 51483 225 51561 271
rect 51607 225 51685 271
rect 51731 225 51809 271
rect 51855 225 51933 271
rect 51979 225 52057 271
rect 52103 225 52181 271
rect 52227 225 52305 271
rect 52351 225 52429 271
rect 52475 225 52553 271
rect 52599 225 52677 271
rect 52723 225 52801 271
rect 52847 225 52925 271
rect 52971 225 53049 271
rect 53095 225 53173 271
rect 53219 225 53297 271
rect 53343 225 53421 271
rect 53467 225 53545 271
rect 53591 225 53669 271
rect 53715 225 53793 271
rect 53839 225 53917 271
rect 53963 225 54041 271
rect 54087 225 54165 271
rect 54211 225 54289 271
rect 54335 225 54413 271
rect 54459 225 54537 271
rect 54583 225 54661 271
rect 54707 225 54785 271
rect 54831 225 54909 271
rect 54955 225 55033 271
rect 55079 225 55157 271
rect 55203 225 55281 271
rect 55327 225 55405 271
rect 55451 225 55529 271
rect 55575 225 55653 271
rect 55699 225 55777 271
rect 55823 225 55901 271
rect 55947 225 56025 271
rect 56071 225 56149 271
rect 56195 225 56273 271
rect 56319 225 56397 271
rect 56443 225 56521 271
rect 56567 225 56645 271
rect 56691 225 56769 271
rect 56815 225 56893 271
rect 56939 225 57017 271
rect 57063 225 57141 271
rect 57187 225 57265 271
rect 57311 225 57389 271
rect 57435 225 57513 271
rect 57559 225 57637 271
rect 57683 225 57761 271
rect 57807 225 57885 271
rect 57931 225 58009 271
rect 58055 225 58133 271
rect 58179 225 58257 271
rect 58303 225 58381 271
rect 58427 225 58505 271
rect 58551 225 58629 271
rect 58675 225 58753 271
rect 58799 225 58877 271
rect 58923 225 59001 271
rect 59047 225 59125 271
rect 59171 225 59249 271
rect 59295 225 59373 271
rect 59419 225 59497 271
rect 59543 225 59621 271
rect 59667 225 59745 271
rect 59791 225 59869 271
rect 59915 225 59993 271
rect 60039 225 60117 271
rect 60163 225 60241 271
rect 60287 225 60365 271
rect 60411 225 60489 271
rect 60535 225 60613 271
rect 60659 225 60737 271
rect 60783 225 60861 271
rect 60907 225 60985 271
rect 61031 225 61109 271
rect 61155 225 61233 271
rect 61279 225 61357 271
rect 61403 225 61481 271
rect 61527 225 61605 271
rect 61651 225 61729 271
rect 61775 225 61853 271
rect 61899 225 61977 271
rect 62023 225 62101 271
rect 62147 225 62225 271
rect 62271 225 62349 271
rect 62395 225 62473 271
rect 62519 225 62597 271
rect 62643 225 62721 271
rect 62767 225 62845 271
rect 62891 225 62969 271
rect 63015 225 63093 271
rect 63139 225 63217 271
rect 63263 225 63341 271
rect 63387 225 63465 271
rect 63511 225 63589 271
rect 63635 225 63713 271
rect 63759 225 63837 271
rect 63883 225 63961 271
rect 64007 225 64085 271
rect 64131 225 64209 271
rect 64255 225 64333 271
rect 64379 225 64457 271
rect 64503 225 64581 271
rect 64627 225 64705 271
rect 64751 225 64829 271
rect 64875 225 64953 271
rect 64999 225 65077 271
rect 65123 225 65201 271
rect 65247 225 65325 271
rect 65371 225 65449 271
rect 65495 225 65573 271
rect 65619 225 65697 271
rect 65743 225 65821 271
rect 65867 225 65945 271
rect 65991 225 66069 271
rect 66115 225 66193 271
rect 66239 225 66317 271
rect 66363 225 66441 271
rect 66487 225 66565 271
rect 66611 225 66689 271
rect 66735 225 66813 271
rect 66859 225 66937 271
rect 66983 225 67061 271
rect 67107 225 67185 271
rect 67231 225 67309 271
rect 67355 225 67433 271
rect 67479 225 67557 271
rect 67603 225 67681 271
rect 67727 225 67805 271
rect 67851 225 67929 271
rect 67975 225 68053 271
rect 68099 225 68177 271
rect 68223 225 68301 271
rect 68347 225 68425 271
rect 68471 225 68549 271
rect 68595 225 68673 271
rect 68719 225 68797 271
rect 68843 225 68921 271
rect 68967 225 69045 271
rect 69091 225 69169 271
rect 69215 225 69293 271
rect 69339 225 69417 271
rect 69463 225 69541 271
rect 69587 225 69665 271
rect 69711 225 69789 271
rect 69835 225 69913 271
rect 69959 225 70037 271
rect 70083 225 70161 271
rect 70207 225 70285 271
rect 70331 225 70409 271
rect 70455 225 70533 271
rect 70579 225 70657 271
rect 70703 225 70781 271
rect 70827 225 70905 271
rect 70951 225 71029 271
rect 71075 225 71153 271
rect 71199 225 71277 271
rect 71323 225 71401 271
rect 71447 225 71525 271
rect 71571 225 71649 271
rect 71695 225 71773 271
rect 71819 225 71897 271
rect 71943 225 72021 271
rect 72067 225 72145 271
rect 72191 225 72269 271
rect 72315 225 72393 271
rect 72439 225 72517 271
rect 72563 225 72641 271
rect 72687 225 72765 271
rect 72811 225 72889 271
rect 72935 225 73013 271
rect 73059 225 73137 271
rect 73183 225 73261 271
rect 73307 225 73385 271
rect 73431 225 73509 271
rect 73555 225 73633 271
rect 73679 225 73757 271
rect 73803 225 73881 271
rect 73927 225 74005 271
rect 74051 225 74129 271
rect 74175 225 74253 271
rect 74299 225 74377 271
rect 74423 225 74501 271
rect 74547 225 74625 271
rect 74671 225 74749 271
rect 74795 225 74873 271
rect 74919 225 74997 271
rect 75043 225 75121 271
rect 75167 225 75245 271
rect 75291 225 75369 271
rect 75415 225 75493 271
rect 75539 225 75617 271
rect 75663 225 75741 271
rect 75787 225 75865 271
rect 75911 225 75989 271
rect 76035 225 76113 271
rect 76159 225 76237 271
rect 76283 225 76361 271
rect 76407 225 76485 271
rect 76531 225 76609 271
rect 76655 225 76733 271
rect 76779 225 76857 271
rect 76903 225 76981 271
rect 77027 225 77105 271
rect 77151 225 77229 271
rect 77275 225 77353 271
rect 77399 225 77477 271
rect 77523 225 77601 271
rect 77647 225 77725 271
rect 77771 225 77849 271
rect 77895 225 77973 271
rect 78019 225 78097 271
rect 78143 225 78221 271
rect 78267 225 78345 271
rect 78391 225 78469 271
rect 78515 225 78593 271
rect 78639 225 78717 271
rect 78763 225 78841 271
rect 78887 225 78965 271
rect 79011 225 79089 271
rect 79135 225 79213 271
rect 79259 225 79337 271
rect 79383 225 79461 271
rect 79507 225 79585 271
rect 79631 225 79709 271
rect 79755 225 79833 271
rect 79879 225 79957 271
rect 80003 225 80081 271
rect 80127 225 80205 271
rect 80251 225 80329 271
rect 80375 225 80453 271
rect 80499 225 80577 271
rect 80623 225 80701 271
rect 80747 225 80825 271
rect 80871 225 80949 271
rect 80995 225 81073 271
rect 81119 225 81197 271
rect 81243 225 81321 271
rect 81367 225 81445 271
rect 81491 225 81569 271
rect 81615 225 81693 271
rect 81739 225 81817 271
rect 81863 225 81941 271
rect 81987 225 82065 271
rect 82111 225 82189 271
rect 82235 225 82313 271
rect 82359 225 82437 271
rect 82483 225 82561 271
rect 82607 225 82685 271
rect 82731 225 82809 271
rect 82855 225 82933 271
rect 82979 225 83057 271
rect 83103 225 83181 271
rect 83227 225 83305 271
rect 83351 225 83429 271
rect 83475 225 83553 271
rect 83599 225 83677 271
rect 83723 225 83801 271
rect 83847 225 83925 271
rect 83971 225 84049 271
rect 84095 225 84173 271
rect 84219 225 84297 271
rect 84343 225 84421 271
rect 84467 225 84545 271
rect 84591 225 84669 271
rect 84715 225 84793 271
rect 84839 225 84917 271
rect 84963 225 85041 271
rect 85087 225 85165 271
rect 85211 225 85289 271
rect 85335 225 85413 271
rect 85459 225 85537 271
rect 85583 225 85594 271
rect -34 147 85594 225
rect -34 101 -23 147
rect 23 101 101 147
rect 147 101 225 147
rect 271 101 349 147
rect 395 101 473 147
rect 519 101 597 147
rect 643 101 721 147
rect 767 101 845 147
rect 891 101 969 147
rect 1015 101 1093 147
rect 1139 101 1217 147
rect 1263 101 1341 147
rect 1387 101 1465 147
rect 1511 101 1589 147
rect 1635 101 1713 147
rect 1759 101 1837 147
rect 1883 101 1961 147
rect 2007 101 2085 147
rect 2131 101 2209 147
rect 2255 101 2333 147
rect 2379 101 2457 147
rect 2503 101 2581 147
rect 2627 101 2705 147
rect 2751 101 2829 147
rect 2875 101 2953 147
rect 2999 101 3077 147
rect 3123 101 3201 147
rect 3247 101 3325 147
rect 3371 101 3449 147
rect 3495 101 3573 147
rect 3619 101 3697 147
rect 3743 101 3821 147
rect 3867 101 3945 147
rect 3991 101 4069 147
rect 4115 101 4193 147
rect 4239 101 4317 147
rect 4363 101 4441 147
rect 4487 101 4565 147
rect 4611 101 4689 147
rect 4735 101 4813 147
rect 4859 101 4937 147
rect 4983 101 5061 147
rect 5107 101 5185 147
rect 5231 101 5309 147
rect 5355 101 5433 147
rect 5479 101 5557 147
rect 5603 101 5681 147
rect 5727 101 5805 147
rect 5851 101 5929 147
rect 5975 101 6053 147
rect 6099 101 6177 147
rect 6223 101 6301 147
rect 6347 101 6425 147
rect 6471 101 6549 147
rect 6595 101 6673 147
rect 6719 101 6797 147
rect 6843 101 6921 147
rect 6967 101 7045 147
rect 7091 101 7169 147
rect 7215 101 7293 147
rect 7339 101 7417 147
rect 7463 101 7541 147
rect 7587 101 7665 147
rect 7711 101 7789 147
rect 7835 101 7913 147
rect 7959 101 8037 147
rect 8083 101 8161 147
rect 8207 101 8285 147
rect 8331 101 8409 147
rect 8455 101 8533 147
rect 8579 101 8657 147
rect 8703 101 8781 147
rect 8827 101 8905 147
rect 8951 101 9029 147
rect 9075 101 9153 147
rect 9199 101 9277 147
rect 9323 101 9401 147
rect 9447 101 9525 147
rect 9571 101 9649 147
rect 9695 101 9773 147
rect 9819 101 9897 147
rect 9943 101 10021 147
rect 10067 101 10145 147
rect 10191 101 10269 147
rect 10315 101 10393 147
rect 10439 101 10517 147
rect 10563 101 10641 147
rect 10687 101 10765 147
rect 10811 101 10889 147
rect 10935 101 11013 147
rect 11059 101 11137 147
rect 11183 101 11261 147
rect 11307 101 11385 147
rect 11431 101 11509 147
rect 11555 101 11633 147
rect 11679 101 11757 147
rect 11803 101 11881 147
rect 11927 101 12005 147
rect 12051 101 12129 147
rect 12175 101 12253 147
rect 12299 101 12377 147
rect 12423 101 12501 147
rect 12547 101 12625 147
rect 12671 101 12749 147
rect 12795 101 12873 147
rect 12919 101 12997 147
rect 13043 101 13121 147
rect 13167 101 13245 147
rect 13291 101 13369 147
rect 13415 101 13493 147
rect 13539 101 13617 147
rect 13663 101 13741 147
rect 13787 101 13865 147
rect 13911 101 13989 147
rect 14035 101 14113 147
rect 14159 101 14237 147
rect 14283 101 14361 147
rect 14407 101 14485 147
rect 14531 101 14609 147
rect 14655 101 14733 147
rect 14779 101 14857 147
rect 14903 101 14981 147
rect 15027 101 15105 147
rect 15151 101 15229 147
rect 15275 101 15353 147
rect 15399 101 15477 147
rect 15523 101 15601 147
rect 15647 101 15725 147
rect 15771 101 15849 147
rect 15895 101 15973 147
rect 16019 101 16097 147
rect 16143 101 16221 147
rect 16267 101 16345 147
rect 16391 101 16469 147
rect 16515 101 16593 147
rect 16639 101 16717 147
rect 16763 101 16841 147
rect 16887 101 16965 147
rect 17011 101 17089 147
rect 17135 101 17213 147
rect 17259 101 17337 147
rect 17383 101 17461 147
rect 17507 101 17585 147
rect 17631 101 17709 147
rect 17755 101 17833 147
rect 17879 101 17957 147
rect 18003 101 18081 147
rect 18127 101 18205 147
rect 18251 101 18329 147
rect 18375 101 18453 147
rect 18499 101 18577 147
rect 18623 101 18701 147
rect 18747 101 18825 147
rect 18871 101 18949 147
rect 18995 101 19073 147
rect 19119 101 19197 147
rect 19243 101 19321 147
rect 19367 101 19445 147
rect 19491 101 19569 147
rect 19615 101 19693 147
rect 19739 101 19817 147
rect 19863 101 19941 147
rect 19987 101 20065 147
rect 20111 101 20189 147
rect 20235 101 20313 147
rect 20359 101 20437 147
rect 20483 101 20561 147
rect 20607 101 20685 147
rect 20731 101 20809 147
rect 20855 101 20933 147
rect 20979 101 21057 147
rect 21103 101 21181 147
rect 21227 101 21305 147
rect 21351 101 21429 147
rect 21475 101 21553 147
rect 21599 101 21677 147
rect 21723 101 21801 147
rect 21847 101 21925 147
rect 21971 101 22049 147
rect 22095 101 22173 147
rect 22219 101 22297 147
rect 22343 101 22421 147
rect 22467 101 22545 147
rect 22591 101 22669 147
rect 22715 101 22793 147
rect 22839 101 22917 147
rect 22963 101 23041 147
rect 23087 101 23165 147
rect 23211 101 23289 147
rect 23335 101 23413 147
rect 23459 101 23537 147
rect 23583 101 23661 147
rect 23707 101 23785 147
rect 23831 101 23909 147
rect 23955 101 24033 147
rect 24079 101 24157 147
rect 24203 101 24281 147
rect 24327 101 24405 147
rect 24451 101 24529 147
rect 24575 101 24653 147
rect 24699 101 24777 147
rect 24823 101 24901 147
rect 24947 101 25025 147
rect 25071 101 25149 147
rect 25195 101 25273 147
rect 25319 101 25397 147
rect 25443 101 25521 147
rect 25567 101 25645 147
rect 25691 101 25769 147
rect 25815 101 25893 147
rect 25939 101 26017 147
rect 26063 101 26141 147
rect 26187 101 26265 147
rect 26311 101 26389 147
rect 26435 101 26513 147
rect 26559 101 26637 147
rect 26683 101 26761 147
rect 26807 101 26885 147
rect 26931 101 27009 147
rect 27055 101 27133 147
rect 27179 101 27257 147
rect 27303 101 27381 147
rect 27427 101 27505 147
rect 27551 101 27629 147
rect 27675 101 27753 147
rect 27799 101 27877 147
rect 27923 101 28001 147
rect 28047 101 28125 147
rect 28171 101 28249 147
rect 28295 101 28373 147
rect 28419 101 28497 147
rect 28543 101 28621 147
rect 28667 101 28745 147
rect 28791 101 28869 147
rect 28915 101 28993 147
rect 29039 101 29117 147
rect 29163 101 29241 147
rect 29287 101 29365 147
rect 29411 101 29489 147
rect 29535 101 29613 147
rect 29659 101 29737 147
rect 29783 101 29861 147
rect 29907 101 29985 147
rect 30031 101 30109 147
rect 30155 101 30233 147
rect 30279 101 30357 147
rect 30403 101 30481 147
rect 30527 101 30605 147
rect 30651 101 30729 147
rect 30775 101 30853 147
rect 30899 101 30977 147
rect 31023 101 31101 147
rect 31147 101 31225 147
rect 31271 101 31349 147
rect 31395 101 31473 147
rect 31519 101 31597 147
rect 31643 101 31721 147
rect 31767 101 31845 147
rect 31891 101 31969 147
rect 32015 101 32093 147
rect 32139 101 32217 147
rect 32263 101 32341 147
rect 32387 101 32465 147
rect 32511 101 32589 147
rect 32635 101 32713 147
rect 32759 101 32837 147
rect 32883 101 32961 147
rect 33007 101 33085 147
rect 33131 101 33209 147
rect 33255 101 33333 147
rect 33379 101 33457 147
rect 33503 101 33581 147
rect 33627 101 33705 147
rect 33751 101 33829 147
rect 33875 101 33953 147
rect 33999 101 34077 147
rect 34123 101 34201 147
rect 34247 101 34325 147
rect 34371 101 34449 147
rect 34495 101 34573 147
rect 34619 101 34697 147
rect 34743 101 34821 147
rect 34867 101 34945 147
rect 34991 101 35069 147
rect 35115 101 35193 147
rect 35239 101 35317 147
rect 35363 101 35441 147
rect 35487 101 35565 147
rect 35611 101 35689 147
rect 35735 101 35813 147
rect 35859 101 35937 147
rect 35983 101 36061 147
rect 36107 101 36185 147
rect 36231 101 36309 147
rect 36355 101 36433 147
rect 36479 101 36557 147
rect 36603 101 36681 147
rect 36727 101 36805 147
rect 36851 101 36929 147
rect 36975 101 37053 147
rect 37099 101 37177 147
rect 37223 101 37301 147
rect 37347 101 37425 147
rect 37471 101 37549 147
rect 37595 101 37673 147
rect 37719 101 37797 147
rect 37843 101 37921 147
rect 37967 101 38045 147
rect 38091 101 38169 147
rect 38215 101 38293 147
rect 38339 101 38417 147
rect 38463 101 38541 147
rect 38587 101 38665 147
rect 38711 101 38789 147
rect 38835 101 38913 147
rect 38959 101 39037 147
rect 39083 101 39161 147
rect 39207 101 39285 147
rect 39331 101 39409 147
rect 39455 101 39533 147
rect 39579 101 39657 147
rect 39703 101 39781 147
rect 39827 101 39905 147
rect 39951 101 40029 147
rect 40075 101 40153 147
rect 40199 101 40277 147
rect 40323 101 40401 147
rect 40447 101 40525 147
rect 40571 101 40649 147
rect 40695 101 40773 147
rect 40819 101 40897 147
rect 40943 101 41021 147
rect 41067 101 41145 147
rect 41191 101 41269 147
rect 41315 101 41393 147
rect 41439 101 41517 147
rect 41563 101 41641 147
rect 41687 101 41765 147
rect 41811 101 41889 147
rect 41935 101 42013 147
rect 42059 101 42137 147
rect 42183 101 42261 147
rect 42307 101 42385 147
rect 42431 101 42509 147
rect 42555 101 42633 147
rect 42679 101 42757 147
rect 42803 101 42881 147
rect 42927 101 43005 147
rect 43051 101 43129 147
rect 43175 101 43253 147
rect 43299 101 43377 147
rect 43423 101 43501 147
rect 43547 101 43625 147
rect 43671 101 43749 147
rect 43795 101 43873 147
rect 43919 101 43997 147
rect 44043 101 44121 147
rect 44167 101 44245 147
rect 44291 101 44369 147
rect 44415 101 44493 147
rect 44539 101 44617 147
rect 44663 101 44741 147
rect 44787 101 44865 147
rect 44911 101 44989 147
rect 45035 101 45113 147
rect 45159 101 45237 147
rect 45283 101 45361 147
rect 45407 101 45485 147
rect 45531 101 45609 147
rect 45655 101 45733 147
rect 45779 101 45857 147
rect 45903 101 45981 147
rect 46027 101 46105 147
rect 46151 101 46229 147
rect 46275 101 46353 147
rect 46399 101 46477 147
rect 46523 101 46601 147
rect 46647 101 46725 147
rect 46771 101 46849 147
rect 46895 101 46973 147
rect 47019 101 47097 147
rect 47143 101 47221 147
rect 47267 101 47345 147
rect 47391 101 47469 147
rect 47515 101 47593 147
rect 47639 101 47717 147
rect 47763 101 47841 147
rect 47887 101 47965 147
rect 48011 101 48089 147
rect 48135 101 48213 147
rect 48259 101 48337 147
rect 48383 101 48461 147
rect 48507 101 48585 147
rect 48631 101 48709 147
rect 48755 101 48833 147
rect 48879 101 48957 147
rect 49003 101 49081 147
rect 49127 101 49205 147
rect 49251 101 49329 147
rect 49375 101 49453 147
rect 49499 101 49577 147
rect 49623 101 49701 147
rect 49747 101 49825 147
rect 49871 101 49949 147
rect 49995 101 50073 147
rect 50119 101 50197 147
rect 50243 101 50321 147
rect 50367 101 50445 147
rect 50491 101 50569 147
rect 50615 101 50693 147
rect 50739 101 50817 147
rect 50863 101 50941 147
rect 50987 101 51065 147
rect 51111 101 51189 147
rect 51235 101 51313 147
rect 51359 101 51437 147
rect 51483 101 51561 147
rect 51607 101 51685 147
rect 51731 101 51809 147
rect 51855 101 51933 147
rect 51979 101 52057 147
rect 52103 101 52181 147
rect 52227 101 52305 147
rect 52351 101 52429 147
rect 52475 101 52553 147
rect 52599 101 52677 147
rect 52723 101 52801 147
rect 52847 101 52925 147
rect 52971 101 53049 147
rect 53095 101 53173 147
rect 53219 101 53297 147
rect 53343 101 53421 147
rect 53467 101 53545 147
rect 53591 101 53669 147
rect 53715 101 53793 147
rect 53839 101 53917 147
rect 53963 101 54041 147
rect 54087 101 54165 147
rect 54211 101 54289 147
rect 54335 101 54413 147
rect 54459 101 54537 147
rect 54583 101 54661 147
rect 54707 101 54785 147
rect 54831 101 54909 147
rect 54955 101 55033 147
rect 55079 101 55157 147
rect 55203 101 55281 147
rect 55327 101 55405 147
rect 55451 101 55529 147
rect 55575 101 55653 147
rect 55699 101 55777 147
rect 55823 101 55901 147
rect 55947 101 56025 147
rect 56071 101 56149 147
rect 56195 101 56273 147
rect 56319 101 56397 147
rect 56443 101 56521 147
rect 56567 101 56645 147
rect 56691 101 56769 147
rect 56815 101 56893 147
rect 56939 101 57017 147
rect 57063 101 57141 147
rect 57187 101 57265 147
rect 57311 101 57389 147
rect 57435 101 57513 147
rect 57559 101 57637 147
rect 57683 101 57761 147
rect 57807 101 57885 147
rect 57931 101 58009 147
rect 58055 101 58133 147
rect 58179 101 58257 147
rect 58303 101 58381 147
rect 58427 101 58505 147
rect 58551 101 58629 147
rect 58675 101 58753 147
rect 58799 101 58877 147
rect 58923 101 59001 147
rect 59047 101 59125 147
rect 59171 101 59249 147
rect 59295 101 59373 147
rect 59419 101 59497 147
rect 59543 101 59621 147
rect 59667 101 59745 147
rect 59791 101 59869 147
rect 59915 101 59993 147
rect 60039 101 60117 147
rect 60163 101 60241 147
rect 60287 101 60365 147
rect 60411 101 60489 147
rect 60535 101 60613 147
rect 60659 101 60737 147
rect 60783 101 60861 147
rect 60907 101 60985 147
rect 61031 101 61109 147
rect 61155 101 61233 147
rect 61279 101 61357 147
rect 61403 101 61481 147
rect 61527 101 61605 147
rect 61651 101 61729 147
rect 61775 101 61853 147
rect 61899 101 61977 147
rect 62023 101 62101 147
rect 62147 101 62225 147
rect 62271 101 62349 147
rect 62395 101 62473 147
rect 62519 101 62597 147
rect 62643 101 62721 147
rect 62767 101 62845 147
rect 62891 101 62969 147
rect 63015 101 63093 147
rect 63139 101 63217 147
rect 63263 101 63341 147
rect 63387 101 63465 147
rect 63511 101 63589 147
rect 63635 101 63713 147
rect 63759 101 63837 147
rect 63883 101 63961 147
rect 64007 101 64085 147
rect 64131 101 64209 147
rect 64255 101 64333 147
rect 64379 101 64457 147
rect 64503 101 64581 147
rect 64627 101 64705 147
rect 64751 101 64829 147
rect 64875 101 64953 147
rect 64999 101 65077 147
rect 65123 101 65201 147
rect 65247 101 65325 147
rect 65371 101 65449 147
rect 65495 101 65573 147
rect 65619 101 65697 147
rect 65743 101 65821 147
rect 65867 101 65945 147
rect 65991 101 66069 147
rect 66115 101 66193 147
rect 66239 101 66317 147
rect 66363 101 66441 147
rect 66487 101 66565 147
rect 66611 101 66689 147
rect 66735 101 66813 147
rect 66859 101 66937 147
rect 66983 101 67061 147
rect 67107 101 67185 147
rect 67231 101 67309 147
rect 67355 101 67433 147
rect 67479 101 67557 147
rect 67603 101 67681 147
rect 67727 101 67805 147
rect 67851 101 67929 147
rect 67975 101 68053 147
rect 68099 101 68177 147
rect 68223 101 68301 147
rect 68347 101 68425 147
rect 68471 101 68549 147
rect 68595 101 68673 147
rect 68719 101 68797 147
rect 68843 101 68921 147
rect 68967 101 69045 147
rect 69091 101 69169 147
rect 69215 101 69293 147
rect 69339 101 69417 147
rect 69463 101 69541 147
rect 69587 101 69665 147
rect 69711 101 69789 147
rect 69835 101 69913 147
rect 69959 101 70037 147
rect 70083 101 70161 147
rect 70207 101 70285 147
rect 70331 101 70409 147
rect 70455 101 70533 147
rect 70579 101 70657 147
rect 70703 101 70781 147
rect 70827 101 70905 147
rect 70951 101 71029 147
rect 71075 101 71153 147
rect 71199 101 71277 147
rect 71323 101 71401 147
rect 71447 101 71525 147
rect 71571 101 71649 147
rect 71695 101 71773 147
rect 71819 101 71897 147
rect 71943 101 72021 147
rect 72067 101 72145 147
rect 72191 101 72269 147
rect 72315 101 72393 147
rect 72439 101 72517 147
rect 72563 101 72641 147
rect 72687 101 72765 147
rect 72811 101 72889 147
rect 72935 101 73013 147
rect 73059 101 73137 147
rect 73183 101 73261 147
rect 73307 101 73385 147
rect 73431 101 73509 147
rect 73555 101 73633 147
rect 73679 101 73757 147
rect 73803 101 73881 147
rect 73927 101 74005 147
rect 74051 101 74129 147
rect 74175 101 74253 147
rect 74299 101 74377 147
rect 74423 101 74501 147
rect 74547 101 74625 147
rect 74671 101 74749 147
rect 74795 101 74873 147
rect 74919 101 74997 147
rect 75043 101 75121 147
rect 75167 101 75245 147
rect 75291 101 75369 147
rect 75415 101 75493 147
rect 75539 101 75617 147
rect 75663 101 75741 147
rect 75787 101 75865 147
rect 75911 101 75989 147
rect 76035 101 76113 147
rect 76159 101 76237 147
rect 76283 101 76361 147
rect 76407 101 76485 147
rect 76531 101 76609 147
rect 76655 101 76733 147
rect 76779 101 76857 147
rect 76903 101 76981 147
rect 77027 101 77105 147
rect 77151 101 77229 147
rect 77275 101 77353 147
rect 77399 101 77477 147
rect 77523 101 77601 147
rect 77647 101 77725 147
rect 77771 101 77849 147
rect 77895 101 77973 147
rect 78019 101 78097 147
rect 78143 101 78221 147
rect 78267 101 78345 147
rect 78391 101 78469 147
rect 78515 101 78593 147
rect 78639 101 78717 147
rect 78763 101 78841 147
rect 78887 101 78965 147
rect 79011 101 79089 147
rect 79135 101 79213 147
rect 79259 101 79337 147
rect 79383 101 79461 147
rect 79507 101 79585 147
rect 79631 101 79709 147
rect 79755 101 79833 147
rect 79879 101 79957 147
rect 80003 101 80081 147
rect 80127 101 80205 147
rect 80251 101 80329 147
rect 80375 101 80453 147
rect 80499 101 80577 147
rect 80623 101 80701 147
rect 80747 101 80825 147
rect 80871 101 80949 147
rect 80995 101 81073 147
rect 81119 101 81197 147
rect 81243 101 81321 147
rect 81367 101 81445 147
rect 81491 101 81569 147
rect 81615 101 81693 147
rect 81739 101 81817 147
rect 81863 101 81941 147
rect 81987 101 82065 147
rect 82111 101 82189 147
rect 82235 101 82313 147
rect 82359 101 82437 147
rect 82483 101 82561 147
rect 82607 101 82685 147
rect 82731 101 82809 147
rect 82855 101 82933 147
rect 82979 101 83057 147
rect 83103 101 83181 147
rect 83227 101 83305 147
rect 83351 101 83429 147
rect 83475 101 83553 147
rect 83599 101 83677 147
rect 83723 101 83801 147
rect 83847 101 83925 147
rect 83971 101 84049 147
rect 84095 101 84173 147
rect 84219 101 84297 147
rect 84343 101 84421 147
rect 84467 101 84545 147
rect 84591 101 84669 147
rect 84715 101 84793 147
rect 84839 101 84917 147
rect 84963 101 85041 147
rect 85087 101 85165 147
rect 85211 101 85289 147
rect 85335 101 85413 147
rect 85459 101 85537 147
rect 85583 101 85594 147
rect -34 23 85594 101
rect -34 -23 -23 23
rect 23 -23 101 23
rect 147 -23 225 23
rect 271 -23 349 23
rect 395 -23 473 23
rect 519 -23 597 23
rect 643 -23 721 23
rect 767 -23 845 23
rect 891 -23 969 23
rect 1015 -23 1093 23
rect 1139 -23 1217 23
rect 1263 -23 1341 23
rect 1387 -23 1465 23
rect 1511 -23 1589 23
rect 1635 -23 1713 23
rect 1759 -23 1837 23
rect 1883 -23 1961 23
rect 2007 -23 2085 23
rect 2131 -23 2209 23
rect 2255 -23 2333 23
rect 2379 -23 2457 23
rect 2503 -23 2581 23
rect 2627 -23 2705 23
rect 2751 -23 2829 23
rect 2875 -23 2953 23
rect 2999 -23 3077 23
rect 3123 -23 3201 23
rect 3247 -23 3325 23
rect 3371 -23 3449 23
rect 3495 -23 3573 23
rect 3619 -23 3697 23
rect 3743 -23 3821 23
rect 3867 -23 3945 23
rect 3991 -23 4069 23
rect 4115 -23 4193 23
rect 4239 -23 4317 23
rect 4363 -23 4441 23
rect 4487 -23 4565 23
rect 4611 -23 4689 23
rect 4735 -23 4813 23
rect 4859 -23 4937 23
rect 4983 -23 5061 23
rect 5107 -23 5185 23
rect 5231 -23 5309 23
rect 5355 -23 5433 23
rect 5479 -23 5557 23
rect 5603 -23 5681 23
rect 5727 -23 5805 23
rect 5851 -23 5929 23
rect 5975 -23 6053 23
rect 6099 -23 6177 23
rect 6223 -23 6301 23
rect 6347 -23 6425 23
rect 6471 -23 6549 23
rect 6595 -23 6673 23
rect 6719 -23 6797 23
rect 6843 -23 6921 23
rect 6967 -23 7045 23
rect 7091 -23 7169 23
rect 7215 -23 7293 23
rect 7339 -23 7417 23
rect 7463 -23 7541 23
rect 7587 -23 7665 23
rect 7711 -23 7789 23
rect 7835 -23 7913 23
rect 7959 -23 8037 23
rect 8083 -23 8161 23
rect 8207 -23 8285 23
rect 8331 -23 8409 23
rect 8455 -23 8533 23
rect 8579 -23 8657 23
rect 8703 -23 8781 23
rect 8827 -23 8905 23
rect 8951 -23 9029 23
rect 9075 -23 9153 23
rect 9199 -23 9277 23
rect 9323 -23 9401 23
rect 9447 -23 9525 23
rect 9571 -23 9649 23
rect 9695 -23 9773 23
rect 9819 -23 9897 23
rect 9943 -23 10021 23
rect 10067 -23 10145 23
rect 10191 -23 10269 23
rect 10315 -23 10393 23
rect 10439 -23 10517 23
rect 10563 -23 10641 23
rect 10687 -23 10765 23
rect 10811 -23 10889 23
rect 10935 -23 11013 23
rect 11059 -23 11137 23
rect 11183 -23 11261 23
rect 11307 -23 11385 23
rect 11431 -23 11509 23
rect 11555 -23 11633 23
rect 11679 -23 11757 23
rect 11803 -23 11881 23
rect 11927 -23 12005 23
rect 12051 -23 12129 23
rect 12175 -23 12253 23
rect 12299 -23 12377 23
rect 12423 -23 12501 23
rect 12547 -23 12625 23
rect 12671 -23 12749 23
rect 12795 -23 12873 23
rect 12919 -23 12997 23
rect 13043 -23 13121 23
rect 13167 -23 13245 23
rect 13291 -23 13369 23
rect 13415 -23 13493 23
rect 13539 -23 13617 23
rect 13663 -23 13741 23
rect 13787 -23 13865 23
rect 13911 -23 13989 23
rect 14035 -23 14113 23
rect 14159 -23 14237 23
rect 14283 -23 14361 23
rect 14407 -23 14485 23
rect 14531 -23 14609 23
rect 14655 -23 14733 23
rect 14779 -23 14857 23
rect 14903 -23 14981 23
rect 15027 -23 15105 23
rect 15151 -23 15229 23
rect 15275 -23 15353 23
rect 15399 -23 15477 23
rect 15523 -23 15601 23
rect 15647 -23 15725 23
rect 15771 -23 15849 23
rect 15895 -23 15973 23
rect 16019 -23 16097 23
rect 16143 -23 16221 23
rect 16267 -23 16345 23
rect 16391 -23 16469 23
rect 16515 -23 16593 23
rect 16639 -23 16717 23
rect 16763 -23 16841 23
rect 16887 -23 16965 23
rect 17011 -23 17089 23
rect 17135 -23 17213 23
rect 17259 -23 17337 23
rect 17383 -23 17461 23
rect 17507 -23 17585 23
rect 17631 -23 17709 23
rect 17755 -23 17833 23
rect 17879 -23 17957 23
rect 18003 -23 18081 23
rect 18127 -23 18205 23
rect 18251 -23 18329 23
rect 18375 -23 18453 23
rect 18499 -23 18577 23
rect 18623 -23 18701 23
rect 18747 -23 18825 23
rect 18871 -23 18949 23
rect 18995 -23 19073 23
rect 19119 -23 19197 23
rect 19243 -23 19321 23
rect 19367 -23 19445 23
rect 19491 -23 19569 23
rect 19615 -23 19693 23
rect 19739 -23 19817 23
rect 19863 -23 19941 23
rect 19987 -23 20065 23
rect 20111 -23 20189 23
rect 20235 -23 20313 23
rect 20359 -23 20437 23
rect 20483 -23 20561 23
rect 20607 -23 20685 23
rect 20731 -23 20809 23
rect 20855 -23 20933 23
rect 20979 -23 21057 23
rect 21103 -23 21181 23
rect 21227 -23 21305 23
rect 21351 -23 21429 23
rect 21475 -23 21553 23
rect 21599 -23 21677 23
rect 21723 -23 21801 23
rect 21847 -23 21925 23
rect 21971 -23 22049 23
rect 22095 -23 22173 23
rect 22219 -23 22297 23
rect 22343 -23 22421 23
rect 22467 -23 22545 23
rect 22591 -23 22669 23
rect 22715 -23 22793 23
rect 22839 -23 22917 23
rect 22963 -23 23041 23
rect 23087 -23 23165 23
rect 23211 -23 23289 23
rect 23335 -23 23413 23
rect 23459 -23 23537 23
rect 23583 -23 23661 23
rect 23707 -23 23785 23
rect 23831 -23 23909 23
rect 23955 -23 24033 23
rect 24079 -23 24157 23
rect 24203 -23 24281 23
rect 24327 -23 24405 23
rect 24451 -23 24529 23
rect 24575 -23 24653 23
rect 24699 -23 24777 23
rect 24823 -23 24901 23
rect 24947 -23 25025 23
rect 25071 -23 25149 23
rect 25195 -23 25273 23
rect 25319 -23 25397 23
rect 25443 -23 25521 23
rect 25567 -23 25645 23
rect 25691 -23 25769 23
rect 25815 -23 25893 23
rect 25939 -23 26017 23
rect 26063 -23 26141 23
rect 26187 -23 26265 23
rect 26311 -23 26389 23
rect 26435 -23 26513 23
rect 26559 -23 26637 23
rect 26683 -23 26761 23
rect 26807 -23 26885 23
rect 26931 -23 27009 23
rect 27055 -23 27133 23
rect 27179 -23 27257 23
rect 27303 -23 27381 23
rect 27427 -23 27505 23
rect 27551 -23 27629 23
rect 27675 -23 27753 23
rect 27799 -23 27877 23
rect 27923 -23 28001 23
rect 28047 -23 28125 23
rect 28171 -23 28249 23
rect 28295 -23 28373 23
rect 28419 -23 28497 23
rect 28543 -23 28621 23
rect 28667 -23 28745 23
rect 28791 -23 28869 23
rect 28915 -23 28993 23
rect 29039 -23 29117 23
rect 29163 -23 29241 23
rect 29287 -23 29365 23
rect 29411 -23 29489 23
rect 29535 -23 29613 23
rect 29659 -23 29737 23
rect 29783 -23 29861 23
rect 29907 -23 29985 23
rect 30031 -23 30109 23
rect 30155 -23 30233 23
rect 30279 -23 30357 23
rect 30403 -23 30481 23
rect 30527 -23 30605 23
rect 30651 -23 30729 23
rect 30775 -23 30853 23
rect 30899 -23 30977 23
rect 31023 -23 31101 23
rect 31147 -23 31225 23
rect 31271 -23 31349 23
rect 31395 -23 31473 23
rect 31519 -23 31597 23
rect 31643 -23 31721 23
rect 31767 -23 31845 23
rect 31891 -23 31969 23
rect 32015 -23 32093 23
rect 32139 -23 32217 23
rect 32263 -23 32341 23
rect 32387 -23 32465 23
rect 32511 -23 32589 23
rect 32635 -23 32713 23
rect 32759 -23 32837 23
rect 32883 -23 32961 23
rect 33007 -23 33085 23
rect 33131 -23 33209 23
rect 33255 -23 33333 23
rect 33379 -23 33457 23
rect 33503 -23 33581 23
rect 33627 -23 33705 23
rect 33751 -23 33829 23
rect 33875 -23 33953 23
rect 33999 -23 34077 23
rect 34123 -23 34201 23
rect 34247 -23 34325 23
rect 34371 -23 34449 23
rect 34495 -23 34573 23
rect 34619 -23 34697 23
rect 34743 -23 34821 23
rect 34867 -23 34945 23
rect 34991 -23 35069 23
rect 35115 -23 35193 23
rect 35239 -23 35317 23
rect 35363 -23 35441 23
rect 35487 -23 35565 23
rect 35611 -23 35689 23
rect 35735 -23 35813 23
rect 35859 -23 35937 23
rect 35983 -23 36061 23
rect 36107 -23 36185 23
rect 36231 -23 36309 23
rect 36355 -23 36433 23
rect 36479 -23 36557 23
rect 36603 -23 36681 23
rect 36727 -23 36805 23
rect 36851 -23 36929 23
rect 36975 -23 37053 23
rect 37099 -23 37177 23
rect 37223 -23 37301 23
rect 37347 -23 37425 23
rect 37471 -23 37549 23
rect 37595 -23 37673 23
rect 37719 -23 37797 23
rect 37843 -23 37921 23
rect 37967 -23 38045 23
rect 38091 -23 38169 23
rect 38215 -23 38293 23
rect 38339 -23 38417 23
rect 38463 -23 38541 23
rect 38587 -23 38665 23
rect 38711 -23 38789 23
rect 38835 -23 38913 23
rect 38959 -23 39037 23
rect 39083 -23 39161 23
rect 39207 -23 39285 23
rect 39331 -23 39409 23
rect 39455 -23 39533 23
rect 39579 -23 39657 23
rect 39703 -23 39781 23
rect 39827 -23 39905 23
rect 39951 -23 40029 23
rect 40075 -23 40153 23
rect 40199 -23 40277 23
rect 40323 -23 40401 23
rect 40447 -23 40525 23
rect 40571 -23 40649 23
rect 40695 -23 40773 23
rect 40819 -23 40897 23
rect 40943 -23 41021 23
rect 41067 -23 41145 23
rect 41191 -23 41269 23
rect 41315 -23 41393 23
rect 41439 -23 41517 23
rect 41563 -23 41641 23
rect 41687 -23 41765 23
rect 41811 -23 41889 23
rect 41935 -23 42013 23
rect 42059 -23 42137 23
rect 42183 -23 42261 23
rect 42307 -23 42385 23
rect 42431 -23 42509 23
rect 42555 -23 42633 23
rect 42679 -23 42757 23
rect 42803 -23 42881 23
rect 42927 -23 43005 23
rect 43051 -23 43129 23
rect 43175 -23 43253 23
rect 43299 -23 43377 23
rect 43423 -23 43501 23
rect 43547 -23 43625 23
rect 43671 -23 43749 23
rect 43795 -23 43873 23
rect 43919 -23 43997 23
rect 44043 -23 44121 23
rect 44167 -23 44245 23
rect 44291 -23 44369 23
rect 44415 -23 44493 23
rect 44539 -23 44617 23
rect 44663 -23 44741 23
rect 44787 -23 44865 23
rect 44911 -23 44989 23
rect 45035 -23 45113 23
rect 45159 -23 45237 23
rect 45283 -23 45361 23
rect 45407 -23 45485 23
rect 45531 -23 45609 23
rect 45655 -23 45733 23
rect 45779 -23 45857 23
rect 45903 -23 45981 23
rect 46027 -23 46105 23
rect 46151 -23 46229 23
rect 46275 -23 46353 23
rect 46399 -23 46477 23
rect 46523 -23 46601 23
rect 46647 -23 46725 23
rect 46771 -23 46849 23
rect 46895 -23 46973 23
rect 47019 -23 47097 23
rect 47143 -23 47221 23
rect 47267 -23 47345 23
rect 47391 -23 47469 23
rect 47515 -23 47593 23
rect 47639 -23 47717 23
rect 47763 -23 47841 23
rect 47887 -23 47965 23
rect 48011 -23 48089 23
rect 48135 -23 48213 23
rect 48259 -23 48337 23
rect 48383 -23 48461 23
rect 48507 -23 48585 23
rect 48631 -23 48709 23
rect 48755 -23 48833 23
rect 48879 -23 48957 23
rect 49003 -23 49081 23
rect 49127 -23 49205 23
rect 49251 -23 49329 23
rect 49375 -23 49453 23
rect 49499 -23 49577 23
rect 49623 -23 49701 23
rect 49747 -23 49825 23
rect 49871 -23 49949 23
rect 49995 -23 50073 23
rect 50119 -23 50197 23
rect 50243 -23 50321 23
rect 50367 -23 50445 23
rect 50491 -23 50569 23
rect 50615 -23 50693 23
rect 50739 -23 50817 23
rect 50863 -23 50941 23
rect 50987 -23 51065 23
rect 51111 -23 51189 23
rect 51235 -23 51313 23
rect 51359 -23 51437 23
rect 51483 -23 51561 23
rect 51607 -23 51685 23
rect 51731 -23 51809 23
rect 51855 -23 51933 23
rect 51979 -23 52057 23
rect 52103 -23 52181 23
rect 52227 -23 52305 23
rect 52351 -23 52429 23
rect 52475 -23 52553 23
rect 52599 -23 52677 23
rect 52723 -23 52801 23
rect 52847 -23 52925 23
rect 52971 -23 53049 23
rect 53095 -23 53173 23
rect 53219 -23 53297 23
rect 53343 -23 53421 23
rect 53467 -23 53545 23
rect 53591 -23 53669 23
rect 53715 -23 53793 23
rect 53839 -23 53917 23
rect 53963 -23 54041 23
rect 54087 -23 54165 23
rect 54211 -23 54289 23
rect 54335 -23 54413 23
rect 54459 -23 54537 23
rect 54583 -23 54661 23
rect 54707 -23 54785 23
rect 54831 -23 54909 23
rect 54955 -23 55033 23
rect 55079 -23 55157 23
rect 55203 -23 55281 23
rect 55327 -23 55405 23
rect 55451 -23 55529 23
rect 55575 -23 55653 23
rect 55699 -23 55777 23
rect 55823 -23 55901 23
rect 55947 -23 56025 23
rect 56071 -23 56149 23
rect 56195 -23 56273 23
rect 56319 -23 56397 23
rect 56443 -23 56521 23
rect 56567 -23 56645 23
rect 56691 -23 56769 23
rect 56815 -23 56893 23
rect 56939 -23 57017 23
rect 57063 -23 57141 23
rect 57187 -23 57265 23
rect 57311 -23 57389 23
rect 57435 -23 57513 23
rect 57559 -23 57637 23
rect 57683 -23 57761 23
rect 57807 -23 57885 23
rect 57931 -23 58009 23
rect 58055 -23 58133 23
rect 58179 -23 58257 23
rect 58303 -23 58381 23
rect 58427 -23 58505 23
rect 58551 -23 58629 23
rect 58675 -23 58753 23
rect 58799 -23 58877 23
rect 58923 -23 59001 23
rect 59047 -23 59125 23
rect 59171 -23 59249 23
rect 59295 -23 59373 23
rect 59419 -23 59497 23
rect 59543 -23 59621 23
rect 59667 -23 59745 23
rect 59791 -23 59869 23
rect 59915 -23 59993 23
rect 60039 -23 60117 23
rect 60163 -23 60241 23
rect 60287 -23 60365 23
rect 60411 -23 60489 23
rect 60535 -23 60613 23
rect 60659 -23 60737 23
rect 60783 -23 60861 23
rect 60907 -23 60985 23
rect 61031 -23 61109 23
rect 61155 -23 61233 23
rect 61279 -23 61357 23
rect 61403 -23 61481 23
rect 61527 -23 61605 23
rect 61651 -23 61729 23
rect 61775 -23 61853 23
rect 61899 -23 61977 23
rect 62023 -23 62101 23
rect 62147 -23 62225 23
rect 62271 -23 62349 23
rect 62395 -23 62473 23
rect 62519 -23 62597 23
rect 62643 -23 62721 23
rect 62767 -23 62845 23
rect 62891 -23 62969 23
rect 63015 -23 63093 23
rect 63139 -23 63217 23
rect 63263 -23 63341 23
rect 63387 -23 63465 23
rect 63511 -23 63589 23
rect 63635 -23 63713 23
rect 63759 -23 63837 23
rect 63883 -23 63961 23
rect 64007 -23 64085 23
rect 64131 -23 64209 23
rect 64255 -23 64333 23
rect 64379 -23 64457 23
rect 64503 -23 64581 23
rect 64627 -23 64705 23
rect 64751 -23 64829 23
rect 64875 -23 64953 23
rect 64999 -23 65077 23
rect 65123 -23 65201 23
rect 65247 -23 65325 23
rect 65371 -23 65449 23
rect 65495 -23 65573 23
rect 65619 -23 65697 23
rect 65743 -23 65821 23
rect 65867 -23 65945 23
rect 65991 -23 66069 23
rect 66115 -23 66193 23
rect 66239 -23 66317 23
rect 66363 -23 66441 23
rect 66487 -23 66565 23
rect 66611 -23 66689 23
rect 66735 -23 66813 23
rect 66859 -23 66937 23
rect 66983 -23 67061 23
rect 67107 -23 67185 23
rect 67231 -23 67309 23
rect 67355 -23 67433 23
rect 67479 -23 67557 23
rect 67603 -23 67681 23
rect 67727 -23 67805 23
rect 67851 -23 67929 23
rect 67975 -23 68053 23
rect 68099 -23 68177 23
rect 68223 -23 68301 23
rect 68347 -23 68425 23
rect 68471 -23 68549 23
rect 68595 -23 68673 23
rect 68719 -23 68797 23
rect 68843 -23 68921 23
rect 68967 -23 69045 23
rect 69091 -23 69169 23
rect 69215 -23 69293 23
rect 69339 -23 69417 23
rect 69463 -23 69541 23
rect 69587 -23 69665 23
rect 69711 -23 69789 23
rect 69835 -23 69913 23
rect 69959 -23 70037 23
rect 70083 -23 70161 23
rect 70207 -23 70285 23
rect 70331 -23 70409 23
rect 70455 -23 70533 23
rect 70579 -23 70657 23
rect 70703 -23 70781 23
rect 70827 -23 70905 23
rect 70951 -23 71029 23
rect 71075 -23 71153 23
rect 71199 -23 71277 23
rect 71323 -23 71401 23
rect 71447 -23 71525 23
rect 71571 -23 71649 23
rect 71695 -23 71773 23
rect 71819 -23 71897 23
rect 71943 -23 72021 23
rect 72067 -23 72145 23
rect 72191 -23 72269 23
rect 72315 -23 72393 23
rect 72439 -23 72517 23
rect 72563 -23 72641 23
rect 72687 -23 72765 23
rect 72811 -23 72889 23
rect 72935 -23 73013 23
rect 73059 -23 73137 23
rect 73183 -23 73261 23
rect 73307 -23 73385 23
rect 73431 -23 73509 23
rect 73555 -23 73633 23
rect 73679 -23 73757 23
rect 73803 -23 73881 23
rect 73927 -23 74005 23
rect 74051 -23 74129 23
rect 74175 -23 74253 23
rect 74299 -23 74377 23
rect 74423 -23 74501 23
rect 74547 -23 74625 23
rect 74671 -23 74749 23
rect 74795 -23 74873 23
rect 74919 -23 74997 23
rect 75043 -23 75121 23
rect 75167 -23 75245 23
rect 75291 -23 75369 23
rect 75415 -23 75493 23
rect 75539 -23 75617 23
rect 75663 -23 75741 23
rect 75787 -23 75865 23
rect 75911 -23 75989 23
rect 76035 -23 76113 23
rect 76159 -23 76237 23
rect 76283 -23 76361 23
rect 76407 -23 76485 23
rect 76531 -23 76609 23
rect 76655 -23 76733 23
rect 76779 -23 76857 23
rect 76903 -23 76981 23
rect 77027 -23 77105 23
rect 77151 -23 77229 23
rect 77275 -23 77353 23
rect 77399 -23 77477 23
rect 77523 -23 77601 23
rect 77647 -23 77725 23
rect 77771 -23 77849 23
rect 77895 -23 77973 23
rect 78019 -23 78097 23
rect 78143 -23 78221 23
rect 78267 -23 78345 23
rect 78391 -23 78469 23
rect 78515 -23 78593 23
rect 78639 -23 78717 23
rect 78763 -23 78841 23
rect 78887 -23 78965 23
rect 79011 -23 79089 23
rect 79135 -23 79213 23
rect 79259 -23 79337 23
rect 79383 -23 79461 23
rect 79507 -23 79585 23
rect 79631 -23 79709 23
rect 79755 -23 79833 23
rect 79879 -23 79957 23
rect 80003 -23 80081 23
rect 80127 -23 80205 23
rect 80251 -23 80329 23
rect 80375 -23 80453 23
rect 80499 -23 80577 23
rect 80623 -23 80701 23
rect 80747 -23 80825 23
rect 80871 -23 80949 23
rect 80995 -23 81073 23
rect 81119 -23 81197 23
rect 81243 -23 81321 23
rect 81367 -23 81445 23
rect 81491 -23 81569 23
rect 81615 -23 81693 23
rect 81739 -23 81817 23
rect 81863 -23 81941 23
rect 81987 -23 82065 23
rect 82111 -23 82189 23
rect 82235 -23 82313 23
rect 82359 -23 82437 23
rect 82483 -23 82561 23
rect 82607 -23 82685 23
rect 82731 -23 82809 23
rect 82855 -23 82933 23
rect 82979 -23 83057 23
rect 83103 -23 83181 23
rect 83227 -23 83305 23
rect 83351 -23 83429 23
rect 83475 -23 83553 23
rect 83599 -23 83677 23
rect 83723 -23 83801 23
rect 83847 -23 83925 23
rect 83971 -23 84049 23
rect 84095 -23 84173 23
rect 84219 -23 84297 23
rect 84343 -23 84421 23
rect 84467 -23 84545 23
rect 84591 -23 84669 23
rect 84715 -23 84793 23
rect 84839 -23 84917 23
rect 84963 -23 85041 23
rect 85087 -23 85165 23
rect 85211 -23 85289 23
rect 85335 -23 85413 23
rect 85459 -23 85537 23
rect 85583 -23 85594 23
rect -34 -34 85594 -23
<< properties >>
string GDS_END 1615338
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1438246
<< end >>
