magic
tech gf180mcuB
timestamp 1667403371
<< metal1 >>
rect 0 111 172 123
rect 11 76 16 104
rect 8 70 18 76
rect 28 70 33 111
rect 11 19 16 70
rect 62 70 67 111
rect 77 70 82 111
rect 133 90 138 111
rect 150 70 160 104
rect 155 64 160 70
rect 155 63 162 64
rect 30 44 40 50
rect 47 43 57 49
rect 49 37 55 43
rect 28 12 33 36
rect 47 31 57 37
rect 154 57 164 63
rect 155 56 162 57
rect 78 44 88 50
rect 104 38 110 48
rect 133 12 138 36
rect 155 19 160 56
rect 0 0 172 12
<< obsm1 >>
rect 45 65 50 104
rect 111 70 121 104
rect 21 59 70 65
rect 111 60 116 70
rect 126 60 136 66
rect 62 19 67 59
rect 94 55 121 60
rect 77 22 82 29
rect 94 27 99 55
rect 115 50 135 55
rect 130 44 145 50
rect 111 22 116 29
rect 77 17 116 22
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 8 69 18 77
rect 154 56 164 64
rect 30 50 40 51
rect 78 50 88 51
rect 30 44 88 50
rect 104 47 110 48
rect 30 43 40 44
rect 78 43 88 44
rect 103 39 111 47
rect 48 37 56 38
rect 103 37 110 39
rect 47 31 110 37
rect 48 30 56 31
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 135 11 143 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 134 5 144 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 135 4 143 5
<< obsm2 >>
rect 60 65 70 66
rect 126 65 136 67
rect 60 59 136 65
rect 60 58 70 59
<< labels >>
rlabel metal2 s 30 43 40 51 6 A
port 1 nsew signal input
rlabel metal2 s 30 44 88 50 6 A
port 1 nsew signal input
rlabel metal2 s 78 43 88 51 6 A
port 1 nsew signal input
rlabel metal1 s 30 44 40 50 6 A
port 1 nsew signal input
rlabel metal1 s 78 44 88 50 6 A
port 1 nsew signal input
rlabel metal2 s 48 30 56 38 6 B
port 2 nsew signal input
rlabel metal2 s 47 31 110 37 6 B
port 2 nsew signal input
rlabel metal2 s 103 31 110 47 6 B
port 2 nsew signal input
rlabel metal2 s 104 31 110 48 6 B
port 2 nsew signal input
rlabel metal2 s 103 39 111 47 6 B
port 2 nsew signal input
rlabel metal1 s 49 31 55 49 6 B
port 2 nsew signal input
rlabel metal1 s 47 31 57 37 6 B
port 2 nsew signal input
rlabel metal1 s 47 43 57 49 6 B
port 2 nsew signal input
rlabel metal1 s 104 38 110 48 6 B
port 2 nsew signal input
rlabel metal2 s 8 69 18 77 6 CO
port 3 nsew signal output
rlabel metal1 s 11 19 16 104 6 CO
port 3 nsew signal output
rlabel metal1 s 8 70 18 76 6 CO
port 3 nsew signal output
rlabel metal2 s 154 56 164 64 6 S
port 4 nsew signal output
rlabel metal1 s 155 19 160 104 6 S
port 4 nsew signal output
rlabel metal1 s 150 70 160 104 6 S
port 4 nsew signal output
rlabel metal1 s 155 56 162 64 6 S
port 4 nsew signal output
rlabel metal1 s 154 57 164 63 6 S
port 4 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 28 70 33 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 62 70 67 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 77 70 82 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 133 90 138 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 111 172 123 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 135 4 143 12 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 134 5 144 11 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 133 0 138 36 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 0 172 12 6 VSS
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 172 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
