magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 5798 870
rect -86 352 2710 377
rect 5447 352 5798 377
<< pwell >>
rect -86 -86 5798 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
rect 1020 68 1140 232
rect 1244 68 1364 232
rect 1468 68 1588 232
rect 1692 68 1812 232
rect 1916 68 2036 232
rect 2140 68 2260 232
rect 2364 68 2484 232
rect 2588 68 2708 232
rect 2916 93 3036 257
rect 3140 93 3260 257
rect 3364 93 3484 257
rect 3588 93 3708 257
rect 3812 93 3932 257
rect 4036 93 4156 257
rect 4260 93 4380 257
rect 4484 93 4604 257
rect 4708 93 4828 257
rect 4932 93 5052 257
rect 5156 93 5276 257
rect 5424 68 5544 232
<< mvpmos >>
rect 144 497 244 716
rect 368 497 468 716
rect 572 497 672 716
rect 816 497 916 716
rect 1020 497 1120 716
rect 1264 497 1364 716
rect 1468 497 1568 716
rect 1692 497 1792 716
rect 1936 497 2036 716
rect 2140 497 2240 716
rect 2384 497 2484 716
rect 2588 497 2688 716
rect 2936 497 3036 716
rect 3140 497 3240 716
rect 3384 497 3484 716
rect 3588 497 3688 716
rect 3832 497 3932 716
rect 4056 497 4156 716
rect 4260 497 4360 716
rect 4504 497 4604 716
rect 4708 497 4808 716
rect 4952 497 5052 716
rect 5156 497 5256 716
rect 5424 497 5524 716
<< mvndiff >>
rect 2816 232 2916 257
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 68 124 173
rect 244 127 348 232
rect 244 81 273 127
rect 319 81 348 127
rect 244 68 348 81
rect 468 219 572 232
rect 468 173 497 219
rect 543 173 572 219
rect 468 68 572 173
rect 692 127 796 232
rect 692 81 721 127
rect 767 81 796 127
rect 692 68 796 81
rect 916 219 1020 232
rect 916 173 945 219
rect 991 173 1020 219
rect 916 68 1020 173
rect 1140 127 1244 232
rect 1140 81 1169 127
rect 1215 81 1244 127
rect 1140 68 1244 81
rect 1364 219 1468 232
rect 1364 173 1393 219
rect 1439 173 1468 219
rect 1364 68 1468 173
rect 1588 127 1692 232
rect 1588 81 1617 127
rect 1663 81 1692 127
rect 1588 68 1692 81
rect 1812 219 1916 232
rect 1812 173 1841 219
rect 1887 173 1916 219
rect 1812 68 1916 173
rect 2036 127 2140 232
rect 2036 81 2065 127
rect 2111 81 2140 127
rect 2036 68 2140 81
rect 2260 219 2364 232
rect 2260 173 2289 219
rect 2335 173 2364 219
rect 2260 68 2364 173
rect 2484 127 2588 232
rect 2484 81 2513 127
rect 2559 81 2588 127
rect 2484 68 2588 81
rect 2708 152 2916 232
rect 2708 106 2747 152
rect 2793 106 2916 152
rect 2708 93 2916 106
rect 3036 244 3140 257
rect 3036 198 3065 244
rect 3111 198 3140 244
rect 3036 93 3140 198
rect 3260 152 3364 257
rect 3260 106 3289 152
rect 3335 106 3364 152
rect 3260 93 3364 106
rect 3484 244 3588 257
rect 3484 198 3513 244
rect 3559 198 3588 244
rect 3484 93 3588 198
rect 3708 152 3812 257
rect 3708 106 3737 152
rect 3783 106 3812 152
rect 3708 93 3812 106
rect 3932 244 4036 257
rect 3932 198 3961 244
rect 4007 198 4036 244
rect 3932 93 4036 198
rect 4156 152 4260 257
rect 4156 106 4185 152
rect 4231 106 4260 152
rect 4156 93 4260 106
rect 4380 244 4484 257
rect 4380 198 4409 244
rect 4455 198 4484 244
rect 4380 93 4484 198
rect 4604 152 4708 257
rect 4604 106 4633 152
rect 4679 106 4708 152
rect 4604 93 4708 106
rect 4828 244 4932 257
rect 4828 198 4857 244
rect 4903 198 4932 244
rect 4828 93 4932 198
rect 5052 152 5156 257
rect 5052 106 5081 152
rect 5127 106 5156 152
rect 5052 93 5156 106
rect 5276 244 5364 257
rect 5276 198 5305 244
rect 5351 232 5364 244
rect 5351 198 5424 232
rect 5276 93 5424 198
rect 2708 68 2808 93
rect 5344 68 5424 93
rect 5544 152 5632 232
rect 5544 106 5573 152
rect 5619 106 5632 152
rect 5544 68 5632 106
<< mvpdiff >>
rect 46 665 144 716
rect 46 525 59 665
rect 105 525 144 665
rect 46 497 144 525
rect 244 497 368 716
rect 468 703 572 716
rect 468 657 497 703
rect 543 657 572 703
rect 468 497 572 657
rect 672 497 816 716
rect 916 664 1020 716
rect 916 618 945 664
rect 991 618 1020 664
rect 916 497 1020 618
rect 1120 497 1264 716
rect 1364 703 1468 716
rect 1364 657 1393 703
rect 1439 657 1468 703
rect 1364 497 1468 657
rect 1568 497 1692 716
rect 1792 497 1936 716
rect 2036 556 2140 716
rect 2036 510 2065 556
rect 2111 510 2140 556
rect 2036 497 2140 510
rect 2240 664 2384 716
rect 2240 618 2289 664
rect 2335 618 2384 664
rect 2240 497 2384 618
rect 2484 556 2588 716
rect 2484 510 2513 556
rect 2559 510 2588 556
rect 2484 497 2588 510
rect 2688 664 2776 716
rect 2688 618 2717 664
rect 2763 618 2776 664
rect 2688 497 2776 618
rect 2848 664 2936 716
rect 2848 618 2861 664
rect 2907 618 2936 664
rect 2848 497 2936 618
rect 3036 556 3140 716
rect 3036 510 3065 556
rect 3111 510 3140 556
rect 3036 497 3140 510
rect 3240 664 3384 716
rect 3240 618 3289 664
rect 3335 618 3384 664
rect 3240 497 3384 618
rect 3484 556 3588 716
rect 3484 510 3513 556
rect 3559 510 3588 556
rect 3484 497 3588 510
rect 3688 497 3832 716
rect 3932 497 4056 716
rect 4156 703 4260 716
rect 4156 657 4185 703
rect 4231 657 4260 703
rect 4156 497 4260 657
rect 4360 497 4504 716
rect 4604 664 4708 716
rect 4604 618 4633 664
rect 4679 618 4708 664
rect 4604 497 4708 618
rect 4808 497 4952 716
rect 5052 703 5156 716
rect 5052 657 5081 703
rect 5127 657 5156 703
rect 5052 497 5156 657
rect 5256 497 5424 716
rect 5524 665 5612 716
rect 5524 525 5553 665
rect 5599 525 5612 665
rect 5524 497 5612 525
<< mvndiffc >>
rect 49 173 95 219
rect 273 81 319 127
rect 497 173 543 219
rect 721 81 767 127
rect 945 173 991 219
rect 1169 81 1215 127
rect 1393 173 1439 219
rect 1617 81 1663 127
rect 1841 173 1887 219
rect 2065 81 2111 127
rect 2289 173 2335 219
rect 2513 81 2559 127
rect 2747 106 2793 152
rect 3065 198 3111 244
rect 3289 106 3335 152
rect 3513 198 3559 244
rect 3737 106 3783 152
rect 3961 198 4007 244
rect 4185 106 4231 152
rect 4409 198 4455 244
rect 4633 106 4679 152
rect 4857 198 4903 244
rect 5081 106 5127 152
rect 5305 198 5351 244
rect 5573 106 5619 152
<< mvpdiffc >>
rect 59 525 105 665
rect 497 657 543 703
rect 945 618 991 664
rect 1393 657 1439 703
rect 2065 510 2111 556
rect 2289 618 2335 664
rect 2513 510 2559 556
rect 2717 618 2763 664
rect 2861 618 2907 664
rect 3065 510 3111 556
rect 3289 618 3335 664
rect 3513 510 3559 556
rect 4185 657 4231 703
rect 4633 618 4679 664
rect 5081 657 5127 703
rect 5553 525 5599 665
<< polysilicon >>
rect 144 716 244 760
rect 368 716 468 760
rect 572 716 672 760
rect 816 716 916 760
rect 1020 716 1120 760
rect 1264 716 1364 760
rect 1468 716 1568 760
rect 1692 716 1792 760
rect 1936 716 2036 760
rect 2140 716 2240 760
rect 2384 716 2484 760
rect 2588 716 2688 760
rect 2936 716 3036 760
rect 3140 716 3240 760
rect 3384 716 3484 760
rect 3588 716 3688 760
rect 3832 716 3932 760
rect 4056 716 4156 760
rect 4260 716 4360 760
rect 4504 716 4604 760
rect 4708 716 4808 760
rect 4952 716 5052 760
rect 5156 716 5256 760
rect 5424 716 5524 760
rect 144 402 244 497
rect 368 415 468 497
rect 368 402 395 415
rect 124 383 244 402
rect 124 337 164 383
rect 210 337 244 383
rect 124 232 244 337
rect 348 369 395 402
rect 441 394 468 415
rect 572 415 672 497
rect 572 394 599 415
rect 441 369 599 394
rect 645 402 672 415
rect 816 433 916 497
rect 816 402 843 433
rect 645 369 692 402
rect 348 348 692 369
rect 348 232 468 348
rect 572 232 692 348
rect 796 387 843 402
rect 889 394 916 433
rect 1020 433 1120 497
rect 1020 394 1047 433
rect 889 387 1047 394
rect 1093 402 1120 433
rect 1264 415 1364 497
rect 1264 402 1291 415
rect 1093 387 1140 402
rect 796 348 1140 387
rect 796 232 916 348
rect 1020 232 1140 348
rect 1244 369 1291 402
rect 1337 394 1364 415
rect 1468 415 1568 497
rect 1468 394 1495 415
rect 1337 369 1495 394
rect 1541 402 1568 415
rect 1692 415 1792 497
rect 1541 369 1588 402
rect 1244 348 1588 369
rect 1244 232 1364 348
rect 1468 232 1588 348
rect 1692 369 1719 415
rect 1765 402 1792 415
rect 1936 415 2036 497
rect 1936 402 1963 415
rect 1765 369 1812 402
rect 1692 232 1812 369
rect 1916 369 1963 402
rect 2009 402 2036 415
rect 2140 415 2240 497
rect 2140 402 2167 415
rect 2009 369 2167 402
rect 2213 402 2240 415
rect 2384 415 2484 497
rect 2384 402 2411 415
rect 2213 369 2411 402
rect 2457 402 2484 415
rect 2588 415 2688 497
rect 2588 402 2608 415
rect 2457 369 2608 402
rect 2654 402 2688 415
rect 2936 415 3036 497
rect 2936 402 2963 415
rect 2654 369 2708 402
rect 1916 348 2708 369
rect 1916 232 2036 348
rect 2140 232 2260 348
rect 2364 232 2484 348
rect 2588 232 2708 348
rect 2916 369 2963 402
rect 3009 402 3036 415
rect 3140 415 3240 497
rect 3140 402 3167 415
rect 3009 369 3167 402
rect 3213 402 3240 415
rect 3384 415 3484 497
rect 3384 402 3411 415
rect 3213 369 3411 402
rect 3457 402 3484 415
rect 3588 415 3688 497
rect 3588 402 3615 415
rect 3457 369 3615 402
rect 3661 402 3688 415
rect 3832 415 3932 497
rect 3832 402 3859 415
rect 3661 369 3708 402
rect 2916 348 3708 369
rect 2916 257 3036 348
rect 3140 257 3260 348
rect 3364 257 3484 348
rect 3588 257 3708 348
rect 3812 369 3859 402
rect 3905 369 3932 415
rect 4056 415 4156 497
rect 4056 402 4083 415
rect 3812 257 3932 369
rect 4036 369 4083 402
rect 4129 394 4156 415
rect 4260 415 4360 497
rect 4260 394 4287 415
rect 4129 369 4287 394
rect 4333 402 4360 415
rect 4504 433 4604 497
rect 4504 402 4531 433
rect 4333 369 4380 402
rect 4036 348 4380 369
rect 4036 257 4156 348
rect 4260 257 4380 348
rect 4484 387 4531 402
rect 4577 394 4604 433
rect 4708 433 4808 497
rect 4708 394 4735 433
rect 4577 387 4735 394
rect 4781 402 4808 433
rect 4952 415 5052 497
rect 4952 402 4979 415
rect 4781 387 4828 402
rect 4484 348 4828 387
rect 4484 257 4604 348
rect 4708 257 4828 348
rect 4932 369 4979 402
rect 5025 394 5052 415
rect 5156 415 5256 497
rect 5156 394 5183 415
rect 5025 369 5183 394
rect 5229 402 5256 415
rect 5424 415 5524 497
rect 5229 369 5276 402
rect 4932 348 5276 369
rect 4932 257 5052 348
rect 5156 257 5276 348
rect 5424 369 5451 415
rect 5497 402 5524 415
rect 5497 369 5544 402
rect 5424 232 5544 369
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
rect 1020 24 1140 68
rect 1244 24 1364 68
rect 1468 24 1588 68
rect 1692 24 1812 68
rect 1916 24 2036 68
rect 2140 24 2260 68
rect 2364 24 2484 68
rect 2588 24 2708 68
rect 2916 24 3036 93
rect 3140 24 3260 93
rect 3364 24 3484 93
rect 3588 24 3708 93
rect 3812 24 3932 93
rect 4036 24 4156 93
rect 4260 24 4380 93
rect 4484 24 4604 93
rect 4708 24 4828 93
rect 4932 24 5052 93
rect 5156 24 5276 93
rect 5424 24 5544 68
<< polycontact >>
rect 164 337 210 383
rect 395 369 441 415
rect 599 369 645 415
rect 843 387 889 433
rect 1047 387 1093 433
rect 1291 369 1337 415
rect 1495 369 1541 415
rect 1719 369 1765 415
rect 1963 369 2009 415
rect 2167 369 2213 415
rect 2411 369 2457 415
rect 2608 369 2654 415
rect 2963 369 3009 415
rect 3167 369 3213 415
rect 3411 369 3457 415
rect 3615 369 3661 415
rect 3859 369 3905 415
rect 4083 369 4129 415
rect 4287 369 4333 415
rect 4531 387 4577 433
rect 4735 387 4781 433
rect 4979 369 5025 415
rect 5183 369 5229 415
rect 5451 369 5497 415
<< metal1 >>
rect 0 724 5712 844
rect 486 703 554 724
rect 59 665 105 676
rect 486 657 497 703
rect 543 657 554 703
rect 1382 703 1450 724
rect 604 618 945 664
rect 991 618 1332 664
rect 1382 657 1393 703
rect 1439 657 1450 703
rect 4174 703 4242 724
rect 604 611 654 618
rect 105 565 654 611
rect 1282 611 1332 618
rect 1500 618 2289 664
rect 2335 618 2717 664
rect 2763 618 2774 664
rect 2848 618 2861 664
rect 2907 618 3289 664
rect 3335 618 4071 664
rect 4174 657 4185 703
rect 4231 657 4242 703
rect 5070 703 5138 724
rect 1500 611 1546 618
rect 1282 565 1546 611
rect 4022 611 4071 618
rect 4292 618 4633 664
rect 4679 618 5020 664
rect 5070 657 5081 703
rect 5127 657 5138 703
rect 5553 665 5599 676
rect 4292 611 4341 618
rect 4022 565 4341 611
rect 4971 611 5020 618
rect 4971 565 5553 611
rect 1916 556 3578 559
rect 59 506 105 525
rect 704 519 1232 540
rect 155 472 1768 519
rect 1916 510 2065 556
rect 2111 510 2513 556
rect 2559 510 3065 556
rect 3111 510 3513 556
rect 3559 510 3578 556
rect 4391 518 4921 542
rect 1916 472 3578 510
rect 3858 472 5498 518
rect 5553 506 5599 525
rect 155 383 219 472
rect 832 433 1104 472
rect 155 337 164 383
rect 210 337 219 383
rect 348 415 764 424
rect 348 369 395 415
rect 441 369 599 415
rect 645 369 764 415
rect 832 387 843 433
rect 889 387 1047 433
rect 1093 387 1104 433
rect 832 384 1104 387
rect 1244 415 1662 424
rect 348 360 764 369
rect 155 306 219 337
rect 718 313 764 360
rect 1244 369 1291 415
rect 1337 369 1495 415
rect 1541 369 1662 415
rect 1244 360 1662 369
rect 1716 415 1768 472
rect 1716 369 1719 415
rect 1765 369 1768 415
rect 1244 313 1290 360
rect 1716 352 1768 369
rect 1916 415 2668 424
rect 1916 369 1963 415
rect 2009 369 2167 415
rect 2213 369 2411 415
rect 2457 369 2608 415
rect 2654 369 2668 415
rect 1916 360 2668 369
rect 718 267 1290 313
rect 2714 244 2774 472
rect 2916 415 3688 424
rect 2916 369 2963 415
rect 3009 369 3167 415
rect 3213 369 3411 415
rect 3457 369 3615 415
rect 3661 369 3688 415
rect 2916 360 3688 369
rect 3858 415 3906 472
rect 4520 433 4792 472
rect 3858 369 3859 415
rect 3905 369 3906 415
rect 3858 352 3906 369
rect 4036 415 4383 424
rect 4036 369 4083 415
rect 4129 369 4287 415
rect 4333 369 4383 415
rect 4520 387 4531 433
rect 4577 387 4735 433
rect 4781 387 4792 433
rect 4520 384 4792 387
rect 4909 415 5367 424
rect 4036 360 4383 369
rect 4337 336 4383 360
rect 4909 369 4979 415
rect 5025 369 5183 415
rect 5229 369 5367 415
rect 4909 360 5367 369
rect 5450 415 5498 472
rect 5450 369 5451 415
rect 5497 369 5498 415
rect 4909 336 4955 360
rect 5450 352 5498 369
rect 4337 290 4955 336
rect 36 173 49 219
rect 95 173 497 219
rect 543 173 945 219
rect 991 173 1393 219
rect 1439 173 1841 219
rect 1887 173 2289 219
rect 2335 173 2666 219
rect 2714 198 3065 244
rect 3111 198 3513 244
rect 3559 198 3961 244
rect 4007 198 4409 244
rect 4455 198 4857 244
rect 4903 198 5305 244
rect 5351 198 5364 244
rect 2620 152 2666 173
rect 262 81 273 127
rect 319 81 330 127
rect 262 60 330 81
rect 710 81 721 127
rect 767 81 778 127
rect 710 60 778 81
rect 1158 81 1169 127
rect 1215 81 1226 127
rect 1158 60 1226 81
rect 1606 81 1617 127
rect 1663 81 1674 127
rect 1606 60 1674 81
rect 2054 81 2065 127
rect 2111 81 2122 127
rect 2054 60 2122 81
rect 2502 81 2513 127
rect 2559 81 2570 127
rect 2620 106 2747 152
rect 2793 106 3289 152
rect 3335 106 3737 152
rect 3783 106 4185 152
rect 4231 106 4633 152
rect 4679 106 5081 152
rect 5127 106 5573 152
rect 5619 106 5632 152
rect 2502 60 2570 81
rect 0 -60 5712 60
<< labels >>
flabel metal1 s 4909 360 5367 424 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 1916 360 2668 424 0 FreeSans 400 0 0 0 B1
port 4 nsew default input
flabel metal1 s 704 519 1232 540 0 FreeSans 400 0 0 0 B2
port 5 nsew default input
flabel metal1 s 1244 360 1662 424 0 FreeSans 400 0 0 0 B3
port 6 nsew default input
flabel metal1 s 0 724 5712 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 2502 60 2570 127 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1916 472 3578 559 0 FreeSans 400 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 2916 360 3688 424 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 4391 518 4921 542 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3858 472 5498 518 1 A2
port 2 nsew default input
rlabel metal1 s 5450 384 5498 472 1 A2
port 2 nsew default input
rlabel metal1 s 4520 384 4792 472 1 A2
port 2 nsew default input
rlabel metal1 s 3858 384 3906 472 1 A2
port 2 nsew default input
rlabel metal1 s 5450 352 5498 384 1 A2
port 2 nsew default input
rlabel metal1 s 3858 352 3906 384 1 A2
port 2 nsew default input
rlabel metal1 s 4036 360 4383 424 1 A3
port 3 nsew default input
rlabel metal1 s 4909 336 4955 360 1 A3
port 3 nsew default input
rlabel metal1 s 4337 336 4383 360 1 A3
port 3 nsew default input
rlabel metal1 s 4337 290 4955 336 1 A3
port 3 nsew default input
rlabel metal1 s 155 472 1768 519 1 B2
port 5 nsew default input
rlabel metal1 s 1716 384 1768 472 1 B2
port 5 nsew default input
rlabel metal1 s 832 384 1104 472 1 B2
port 5 nsew default input
rlabel metal1 s 155 384 219 472 1 B2
port 5 nsew default input
rlabel metal1 s 1716 352 1768 384 1 B2
port 5 nsew default input
rlabel metal1 s 155 352 219 384 1 B2
port 5 nsew default input
rlabel metal1 s 155 306 219 352 1 B2
port 5 nsew default input
rlabel metal1 s 348 360 764 424 1 B3
port 6 nsew default input
rlabel metal1 s 1244 313 1290 360 1 B3
port 6 nsew default input
rlabel metal1 s 718 313 764 360 1 B3
port 6 nsew default input
rlabel metal1 s 718 267 1290 313 1 B3
port 6 nsew default input
rlabel metal1 s 2714 244 2774 472 1 ZN
port 7 nsew default output
rlabel metal1 s 2714 198 5364 244 1 ZN
port 7 nsew default output
rlabel metal1 s 5070 657 5138 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4174 657 4242 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1382 657 1450 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 486 657 554 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2054 60 2122 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1606 60 1674 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1158 60 1226 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 710 60 778 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5712 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5712 784
string GDS_END 87094
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 77580
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
