magic
tech gf180mcuB
timestamp 1667403374
<< metal1 >>
rect 0 147 300 159
rect 11 106 16 147
rect 28 91 33 140
rect 45 106 50 147
rect 62 91 67 140
rect 79 106 84 147
rect 96 91 101 140
rect 113 106 118 147
rect 130 91 135 140
rect 147 106 152 147
rect 164 91 169 140
rect 181 106 186 147
rect 198 91 203 140
rect 215 106 220 147
rect 232 91 237 140
rect 249 106 254 147
rect 266 91 271 140
rect 283 106 288 147
rect 28 86 271 91
rect 8 67 18 73
rect 28 43 33 86
rect 62 43 67 86
rect 96 43 101 86
rect 130 43 135 86
rect 164 43 169 86
rect 198 43 203 86
rect 232 43 237 86
rect 263 84 271 86
rect 266 43 271 84
rect 28 38 271 43
rect 11 9 16 33
rect 28 16 33 38
rect 45 9 50 33
rect 62 16 67 38
rect 79 9 84 33
rect 96 16 101 38
rect 113 9 118 33
rect 130 16 135 38
rect 147 9 152 33
rect 164 16 169 38
rect 181 9 186 33
rect 198 16 203 38
rect 215 9 220 33
rect 232 16 237 38
rect 249 9 254 33
rect 266 16 271 38
rect 283 9 288 33
rect 0 -3 300 9
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 130 154 138 155
rect 154 154 162 155
rect 178 154 186 155
rect 202 154 210 155
rect 226 154 234 155
rect 250 154 258 155
rect 274 154 282 155
rect 9 148 19 154
rect 33 148 43 154
rect 57 148 67 154
rect 81 148 91 154
rect 105 148 115 154
rect 129 148 139 154
rect 153 148 163 154
rect 177 148 187 154
rect 201 148 211 154
rect 225 148 235 154
rect 249 148 259 154
rect 273 148 283 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 130 147 138 148
rect 154 147 162 148
rect 178 147 186 148
rect 202 147 210 148
rect 226 147 234 148
rect 250 147 258 148
rect 274 147 282 148
rect 263 84 273 92
rect 8 66 18 74
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 82 8 90 9
rect 106 8 114 9
rect 130 8 138 9
rect 154 8 162 9
rect 178 8 186 9
rect 202 8 210 9
rect 226 8 234 9
rect 250 8 258 9
rect 274 8 282 9
rect 9 2 19 8
rect 33 2 43 8
rect 57 2 67 8
rect 81 2 91 8
rect 105 2 115 8
rect 129 2 139 8
rect 153 2 163 8
rect 177 2 187 8
rect 201 2 211 8
rect 225 2 235 8
rect 249 2 259 8
rect 273 2 283 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
rect 82 1 90 2
rect 106 1 114 2
rect 130 1 138 2
rect 154 1 162 2
rect 178 1 186 2
rect 202 1 210 2
rect 226 1 234 2
rect 250 1 258 2
rect 274 1 282 2
<< labels >>
rlabel metal2 s 8 66 18 74 6 A
port 1 nsew signal input
rlabel metal1 s 8 67 18 73 6 A
port 1 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 34 147 42 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 33 148 43 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 58 147 66 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 57 148 67 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 82 147 90 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 81 148 91 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 106 147 114 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 105 148 115 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 130 147 138 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 129 148 139 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 154 147 162 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 153 148 163 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 178 147 186 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 177 148 187 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 202 147 210 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 201 148 211 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 226 147 234 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 225 148 235 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 250 147 258 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 249 148 259 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 274 147 282 155 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 273 148 283 154 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 45 106 50 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 79 106 84 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 113 106 118 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 147 106 152 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 181 106 186 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 215 106 220 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 249 106 254 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 283 106 288 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 147 300 159 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 34 1 42 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 33 2 43 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 58 1 66 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 57 2 67 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 82 1 90 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 81 2 91 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 106 1 114 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 105 2 115 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 130 1 138 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 129 2 139 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 154 1 162 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 153 2 163 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 178 1 186 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 177 2 187 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 202 1 210 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 201 2 211 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 226 1 234 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 225 2 235 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 250 1 258 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 249 2 259 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 274 1 282 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 273 2 283 8 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 45 -3 50 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 79 -3 84 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 113 -3 118 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 147 -3 152 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 181 -3 186 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 215 -3 220 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 249 -3 254 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 283 -3 288 33 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 0 -3 300 9 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 263 84 273 92 6 Y
port 4 nsew signal output
rlabel metal1 s 28 16 33 140 6 Y
port 4 nsew signal output
rlabel metal1 s 62 16 67 140 6 Y
port 4 nsew signal output
rlabel metal1 s 96 16 101 140 6 Y
port 4 nsew signal output
rlabel metal1 s 130 16 135 140 6 Y
port 4 nsew signal output
rlabel metal1 s 164 16 169 140 6 Y
port 4 nsew signal output
rlabel metal1 s 198 16 203 140 6 Y
port 4 nsew signal output
rlabel metal1 s 232 16 237 140 6 Y
port 4 nsew signal output
rlabel metal1 s 28 38 271 43 6 Y
port 4 nsew signal output
rlabel metal1 s 263 84 271 91 6 Y
port 4 nsew signal output
rlabel metal1 s 28 86 271 91 6 Y
port 4 nsew signal output
rlabel metal1 s 266 16 271 140 6 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 300 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
