magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 95023 342 95042
rect -42 -23 -23 95023
rect 323 -23 342 95023
rect -42 -42 342 -23
<< psubdiffcont >>
rect -23 -23 323 95023
<< metal1 >>
rect -34 95023 334 95034
rect -34 -23 -23 95023
rect 323 -23 334 95023
rect -34 -34 334 -23
<< properties >>
string GDS_END 1557694
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1314042
<< end >>
