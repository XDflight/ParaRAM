magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 2272 33837 2372 34659
rect 7620 34632 7696 34644
rect 7620 34268 7632 34632
rect 7684 34268 7696 34632
rect 7620 34256 7696 34268
rect 13072 33837 13282 34659
rect 18400 34632 18516 34659
rect 18400 34268 18432 34632
rect 18484 34268 18516 34632
rect 18400 33981 18516 34268
rect 23512 33837 23612 34659
rect 61740 33837 61948 34659
rect 67176 34632 67292 34659
rect 67176 34268 67208 34632
rect 67260 34268 67292 34632
rect 67176 33981 67292 34268
rect 72648 33763 72858 34659
rect 77879 34632 78084 34659
rect 77879 34268 78008 34632
rect 78060 34268 78084 34632
rect 77879 33811 78084 34268
rect 83088 34005 83188 34659
rect 82716 33722 83188 34005
<< via1 >>
rect 7632 34268 7684 34632
rect 18432 34268 18484 34632
rect 67208 34268 67260 34632
rect 78008 34268 78060 34632
<< metal2 >>
rect 7672 35034 7772 35222
rect 18472 35034 18572 35222
rect 67248 35034 67348 35222
rect 78048 35034 78148 35222
rect 7608 34934 7772 35034
rect 18408 34934 18572 35034
rect 67184 34934 67348 35034
rect 77984 34934 78148 35034
rect 7608 34632 7708 34934
rect 7608 34268 7632 34632
rect 7684 34268 7708 34632
rect 7608 34245 7708 34268
rect 18408 34632 18508 34934
rect 18408 34268 18432 34632
rect 18484 34268 18508 34632
rect 18408 34245 18508 34268
rect 1912 26265 2012 32592
rect 12712 32366 12812 32592
rect 12712 32266 13049 32366
rect 12955 31889 13049 32266
rect 23872 31965 23972 32592
rect 23755 31865 23972 31965
rect 12571 28377 12647 28387
rect 12571 28321 12581 28377
rect 12637 28321 12647 28377
rect 12571 28265 12647 28321
rect 12571 28209 12581 28265
rect 12637 28209 12647 28265
rect 12571 28153 12647 28209
rect 12571 28097 12581 28153
rect 12637 28097 12647 28153
rect 12571 28041 12647 28097
rect 12571 27985 12581 28041
rect 12637 27985 12647 28041
rect 12571 27929 12647 27985
rect 12571 27873 12581 27929
rect 12637 27873 12647 27929
rect 12571 27817 12647 27873
rect 12571 27761 12581 27817
rect 12637 27761 12647 27817
rect 12571 27751 12647 27761
rect 12964 28377 13040 28387
rect 12964 28321 12974 28377
rect 13030 28321 13040 28377
rect 12964 28265 13040 28321
rect 12964 28209 12974 28265
rect 13030 28209 13040 28265
rect 12964 28153 13040 28209
rect 12964 28097 12974 28153
rect 13030 28097 13040 28153
rect 12964 28041 13040 28097
rect 12964 27985 12974 28041
rect 13030 27985 13040 28041
rect 12964 27929 13040 27985
rect 12964 27873 12974 27929
rect 13030 27873 13040 27929
rect 12964 27817 13040 27873
rect 12964 27761 12974 27817
rect 13030 27761 13040 27817
rect 12964 27751 13040 27761
rect 23371 28377 23447 28387
rect 23371 28321 23381 28377
rect 23437 28321 23447 28377
rect 23371 28265 23447 28321
rect 23371 28209 23381 28265
rect 23437 28209 23447 28265
rect 23371 28153 23447 28209
rect 23371 28097 23381 28153
rect 23437 28097 23447 28153
rect 23371 28041 23447 28097
rect 23371 27985 23381 28041
rect 23437 27985 23447 28041
rect 23371 27929 23447 27985
rect 23371 27873 23381 27929
rect 23437 27873 23447 27929
rect 23371 27817 23447 27873
rect 23371 27761 23381 27817
rect 23437 27761 23447 27817
rect 23371 27751 23447 27761
rect 23764 28377 23840 28387
rect 23764 28321 23774 28377
rect 23830 28321 23840 28377
rect 23764 28265 23840 28321
rect 23764 28209 23774 28265
rect 23830 28209 23840 28265
rect 23764 28153 23840 28209
rect 23764 28097 23774 28153
rect 23830 28097 23840 28153
rect 23764 28041 23840 28097
rect 23764 27985 23774 28041
rect 23830 27985 23840 28041
rect 23764 27929 23840 27985
rect 23764 27873 23774 27929
rect 23830 27873 23840 27929
rect 23764 27817 23840 27873
rect 23764 27761 23774 27817
rect 23830 27761 23840 27817
rect 23764 27751 23840 27761
rect 61487 26265 61587 34760
rect 67184 34632 67284 34934
rect 67184 34268 67208 34632
rect 67260 34268 67284 34632
rect 67184 34245 67284 34268
rect 72288 32366 72388 34758
rect 77984 34632 78084 34934
rect 77984 34268 78008 34632
rect 78060 34268 78084 34632
rect 77984 34245 78084 34268
rect 72288 32266 72625 32366
rect 72531 31889 72625 32266
rect 83448 31965 83548 32592
rect 83331 31865 83548 31965
rect 72147 28377 72223 28387
rect 72147 28321 72157 28377
rect 72213 28321 72223 28377
rect 72147 28265 72223 28321
rect 72147 28209 72157 28265
rect 72213 28209 72223 28265
rect 72147 28153 72223 28209
rect 72147 28097 72157 28153
rect 72213 28097 72223 28153
rect 72147 28041 72223 28097
rect 72147 27985 72157 28041
rect 72213 27985 72223 28041
rect 72147 27929 72223 27985
rect 72147 27873 72157 27929
rect 72213 27873 72223 27929
rect 72147 27817 72223 27873
rect 72147 27761 72157 27817
rect 72213 27761 72223 27817
rect 72147 27751 72223 27761
rect 72540 28377 72616 28387
rect 72540 28321 72550 28377
rect 72606 28321 72616 28377
rect 72540 28265 72616 28321
rect 72540 28209 72550 28265
rect 72606 28209 72616 28265
rect 72540 28153 72616 28209
rect 72540 28097 72550 28153
rect 72606 28097 72616 28153
rect 72540 28041 72616 28097
rect 72540 27985 72550 28041
rect 72606 27985 72616 28041
rect 72540 27929 72616 27985
rect 72540 27873 72550 27929
rect 72606 27873 72616 27929
rect 72540 27817 72616 27873
rect 72540 27761 72550 27817
rect 72606 27761 72616 27817
rect 72540 27751 72616 27761
rect 82947 28377 83023 28387
rect 82947 28321 82957 28377
rect 83013 28321 83023 28377
rect 82947 28265 83023 28321
rect 82947 28209 82957 28265
rect 83013 28209 83023 28265
rect 82947 28153 83023 28209
rect 82947 28097 82957 28153
rect 83013 28097 83023 28153
rect 82947 28041 83023 28097
rect 82947 27985 82957 28041
rect 83013 27985 83023 28041
rect 82947 27929 83023 27985
rect 82947 27873 82957 27929
rect 83013 27873 83023 27929
rect 82947 27817 83023 27873
rect 82947 27761 82957 27817
rect 83013 27761 83023 27817
rect 82947 27751 83023 27761
rect 83340 28377 83416 28387
rect 83340 28321 83350 28377
rect 83406 28321 83416 28377
rect 83340 28265 83416 28321
rect 83340 28209 83350 28265
rect 83406 28209 83416 28265
rect 83340 28153 83416 28209
rect 83340 28097 83350 28153
rect 83406 28097 83416 28153
rect 83340 28041 83416 28097
rect 83340 27985 83350 28041
rect 83406 27985 83416 28041
rect 83340 27929 83416 27985
rect 83340 27873 83350 27929
rect 83406 27873 83416 27929
rect 83340 27817 83416 27873
rect 83340 27761 83350 27817
rect 83406 27761 83416 27817
rect 83340 27751 83416 27761
<< via2 >>
rect 12581 28321 12637 28377
rect 12581 28209 12637 28265
rect 12581 28097 12637 28153
rect 12581 27985 12637 28041
rect 12581 27873 12637 27929
rect 12581 27761 12637 27817
rect 12974 28321 13030 28377
rect 12974 28209 13030 28265
rect 12974 28097 13030 28153
rect 12974 27985 13030 28041
rect 12974 27873 13030 27929
rect 12974 27761 13030 27817
rect 23381 28321 23437 28377
rect 23381 28209 23437 28265
rect 23381 28097 23437 28153
rect 23381 27985 23437 28041
rect 23381 27873 23437 27929
rect 23381 27761 23437 27817
rect 23774 28321 23830 28377
rect 23774 28209 23830 28265
rect 23774 28097 23830 28153
rect 23774 27985 23830 28041
rect 23774 27873 23830 27929
rect 23774 27761 23830 27817
rect 72157 28321 72213 28377
rect 72157 28209 72213 28265
rect 72157 28097 72213 28153
rect 72157 27985 72213 28041
rect 72157 27873 72213 27929
rect 72157 27761 72213 27817
rect 72550 28321 72606 28377
rect 72550 28209 72606 28265
rect 72550 28097 72606 28153
rect 72550 27985 72606 28041
rect 72550 27873 72606 27929
rect 72550 27761 72606 27817
rect 82957 28321 83013 28377
rect 82957 28209 83013 28265
rect 82957 28097 83013 28153
rect 82957 27985 83013 28041
rect 82957 27873 83013 27929
rect 82957 27761 83013 27817
rect 83350 28321 83406 28377
rect 83350 28209 83406 28265
rect 83350 28097 83406 28153
rect 83350 27985 83406 28041
rect 83350 27873 83406 27929
rect 83350 27761 83406 27817
<< metal3 >>
rect 12571 28377 12647 28387
rect 12571 28321 12581 28377
rect 12637 28321 12647 28377
rect 12571 28265 12647 28321
rect 12571 28209 12581 28265
rect 12637 28209 12647 28265
rect 12571 28153 12647 28209
rect 12571 28097 12581 28153
rect 12637 28097 12647 28153
rect 12571 28041 12647 28097
rect 12571 27985 12581 28041
rect 12637 27985 12647 28041
rect 12571 27929 12647 27985
rect 12571 27873 12581 27929
rect 12637 27873 12647 27929
rect 12571 27817 12647 27873
rect 12571 27761 12581 27817
rect 12637 27761 12647 27817
rect 12571 27751 12647 27761
rect 12964 28377 13040 28387
rect 12964 28321 12974 28377
rect 13030 28321 13040 28377
rect 12964 28265 13040 28321
rect 12964 28209 12974 28265
rect 13030 28209 13040 28265
rect 12964 28153 13040 28209
rect 12964 28097 12974 28153
rect 13030 28097 13040 28153
rect 12964 28041 13040 28097
rect 12964 27985 12974 28041
rect 13030 27985 13040 28041
rect 12964 27929 13040 27985
rect 12964 27873 12974 27929
rect 13030 27873 13040 27929
rect 12964 27817 13040 27873
rect 12964 27761 12974 27817
rect 13030 27761 13040 27817
rect 12964 27751 13040 27761
rect 23371 28377 23447 28387
rect 23371 28321 23381 28377
rect 23437 28321 23447 28377
rect 23371 28265 23447 28321
rect 23371 28209 23381 28265
rect 23437 28209 23447 28265
rect 23371 28153 23447 28209
rect 23371 28097 23381 28153
rect 23437 28097 23447 28153
rect 23371 28041 23447 28097
rect 23371 27985 23381 28041
rect 23437 27985 23447 28041
rect 23371 27929 23447 27985
rect 23371 27873 23381 27929
rect 23437 27873 23447 27929
rect 23371 27817 23447 27873
rect 23371 27761 23381 27817
rect 23437 27761 23447 27817
rect 23371 27751 23447 27761
rect 23764 28377 23840 28387
rect 23764 28321 23774 28377
rect 23830 28321 23840 28377
rect 23764 28265 23840 28321
rect 23764 28209 23774 28265
rect 23830 28209 23840 28265
rect 23764 28153 23840 28209
rect 23764 28097 23774 28153
rect 23830 28097 23840 28153
rect 23764 28041 23840 28097
rect 23764 27985 23774 28041
rect 23830 27985 23840 28041
rect 23764 27929 23840 27985
rect 23764 27873 23774 27929
rect 23830 27873 23840 27929
rect 23764 27817 23840 27873
rect 23764 27761 23774 27817
rect 23830 27761 23840 27817
rect 23764 27751 23840 27761
rect 72147 28377 72223 28387
rect 72147 28321 72157 28377
rect 72213 28321 72223 28377
rect 72147 28265 72223 28321
rect 72147 28209 72157 28265
rect 72213 28209 72223 28265
rect 72147 28153 72223 28209
rect 72147 28097 72157 28153
rect 72213 28097 72223 28153
rect 72147 28041 72223 28097
rect 72147 27985 72157 28041
rect 72213 27985 72223 28041
rect 72147 27929 72223 27985
rect 72147 27873 72157 27929
rect 72213 27873 72223 27929
rect 72147 27817 72223 27873
rect 72147 27761 72157 27817
rect 72213 27761 72223 27817
rect 72147 27751 72223 27761
rect 72540 28377 72616 28387
rect 72540 28321 72550 28377
rect 72606 28321 72616 28377
rect 72540 28265 72616 28321
rect 72540 28209 72550 28265
rect 72606 28209 72616 28265
rect 72540 28153 72616 28209
rect 72540 28097 72550 28153
rect 72606 28097 72616 28153
rect 72540 28041 72616 28097
rect 72540 27985 72550 28041
rect 72606 27985 72616 28041
rect 72540 27929 72616 27985
rect 72540 27873 72550 27929
rect 72606 27873 72616 27929
rect 72540 27817 72616 27873
rect 72540 27761 72550 27817
rect 72606 27761 72616 27817
rect 72540 27751 72616 27761
rect 82947 28377 83023 28387
rect 82947 28321 82957 28377
rect 83013 28321 83023 28377
rect 82947 28265 83023 28321
rect 82947 28209 82957 28265
rect 83013 28209 83023 28265
rect 82947 28153 83023 28209
rect 82947 28097 82957 28153
rect 83013 28097 83023 28153
rect 82947 28041 83023 28097
rect 82947 27985 82957 28041
rect 83013 27985 83023 28041
rect 82947 27929 83023 27985
rect 82947 27873 82957 27929
rect 83013 27873 83023 27929
rect 82947 27817 83023 27873
rect 82947 27761 82957 27817
rect 83013 27761 83023 27817
rect 82947 27751 83023 27761
rect 83340 28377 83416 28387
rect 83340 28321 83350 28377
rect 83406 28321 83416 28377
rect 83340 28265 83416 28321
rect 83340 28209 83350 28265
rect 83406 28209 83416 28265
rect 83340 28153 83416 28209
rect 83340 28097 83350 28153
rect 83406 28097 83416 28153
rect 83340 28041 83416 28097
rect 83340 27985 83350 28041
rect 83406 27985 83416 28041
rect 83340 27929 83416 27985
rect 83340 27873 83350 27929
rect 83406 27873 83416 27929
rect 83340 27817 83416 27873
rect 83340 27761 83350 27817
rect 83406 27761 83416 27817
rect 83340 27751 83416 27761
rect 46982 15015 47947 16784
rect 27546 14936 47947 15015
rect 27546 14503 47683 14936
rect 41493 14491 47683 14503
rect 41493 13729 45977 14491
rect 41151 6592 51232 7392
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_0
timestamp 1666464484
transform 1 0 18458 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_1
timestamp 1666464484
transform 1 0 67234 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_2
timestamp 1666464484
transform 1 0 78034 0 1 34450
box 0 0 1 1
use M2_M14310590878121_256x8m81  M2_M14310590878121_256x8m81_3
timestamp 1666464484
transform 1 0 7658 0 1 34450
box 0 0 1 1
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_0
timestamp 1666464484
transform -1 0 72698 0 1 34224
box -38 -402 38 402
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_1
timestamp 1666464484
transform -1 0 83138 0 1 34224
box -38 -402 38 402
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_2
timestamp 1666464484
transform -1 0 61898 0 1 34224
box -38 -402 38 402
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_3
timestamp 1666464484
transform 1 0 13122 0 1 34224
box -38 -402 38 402
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_4
timestamp 1666464484
transform 1 0 2322 0 1 34224
box -38 -402 38 402
use M2_M14310590878199_256x8m81  M2_M14310590878199_256x8m81_5
timestamp 1666464484
transform 1 0 23562 0 1 34224
box -38 -402 38 402
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_0
timestamp 1666464484
transform 1 0 12609 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_1
timestamp 1666464484
transform 1 0 23802 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_2
timestamp 1666464484
transform 1 0 23409 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_3
timestamp 1666464484
transform 1 0 72578 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_4
timestamp 1666464484
transform 1 0 72185 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_5
timestamp 1666464484
transform 1 0 83378 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_6
timestamp 1666464484
transform 1 0 82985 0 1 26882
box -38 -430 38 430
use M3_M243105908781100_256x8m81  M3_M243105908781100_256x8m81_7
timestamp 1666464484
transform 1 0 13002 0 1 26882
box -38 -430 38 430
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_0
timestamp 1666464484
transform 1 0 12609 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_1
timestamp 1666464484
transform 1 0 23802 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_2
timestamp 1666464484
transform 1 0 23409 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_3
timestamp 1666464484
transform 1 0 72578 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_4
timestamp 1666464484
transform 1 0 72185 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_5
timestamp 1666464484
transform 1 0 83378 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_6
timestamp 1666464484
transform 1 0 82985 0 1 28069
box 0 0 1 1
use M3_M243105908781101_256x8m81  M3_M243105908781101_256x8m81_7
timestamp 1666464484
transform 1 0 13002 0 1 28069
box 0 0 1 1
use M3_M243105908781102_256x8m81  M3_M243105908781102_256x8m81_0
timestamp 1666464484
transform 1 0 61537 0 1 27432
box -38 -908 38 908
use M3_M243105908781102_256x8m81  M3_M243105908781102_256x8m81_1
timestamp 1666464484
transform 1 0 1962 0 1 27432
box -38 -908 38 908
<< properties >>
string GDS_END 2289314
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2286308
string path 205.755 34.960 256.160 34.960 
<< end >>
