magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -143 76 143 81
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -81 143 -76
<< via2 >>
rect -138 48 -110 76
rect -76 48 -48 76
rect -14 48 14 76
rect 48 48 76 76
rect 110 48 138 76
rect -138 -14 -110 14
rect -76 -14 -48 14
rect -14 -14 14 14
rect 48 -14 76 14
rect 110 -14 138 14
rect -138 -76 -110 -48
rect -76 -76 -48 -48
rect -14 -76 14 -48
rect 48 -76 76 -48
rect 110 -76 138 -48
<< metal3 >>
rect -143 76 143 81
rect -143 48 -138 76
rect -110 48 -76 76
rect -48 48 -14 76
rect 14 48 48 76
rect 76 48 110 76
rect 138 48 143 76
rect -143 14 143 48
rect -143 -14 -138 14
rect -110 -14 -76 14
rect -48 -14 -14 14
rect 14 -14 48 14
rect 76 -14 110 14
rect 138 -14 143 14
rect -143 -48 143 -14
rect -143 -76 -138 -48
rect -110 -76 -76 -48
rect -48 -76 -14 -48
rect 14 -76 48 -48
rect 76 -76 110 -48
rect 138 -76 143 -48
rect -143 -81 143 -76
<< properties >>
string GDS_END 1736090
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1734998
<< end >>
