magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 18619 16077 18786 16532
rect 278 4553 5772 7557
rect 458 1191 5467 2381
rect 7020 126 8322 862
<< pmos >>
rect 7275 267 7395 722
rect 7499 267 7619 722
rect 7723 267 7843 722
rect 7947 267 8067 722
<< ndiff >>
rect 18553 16224 18619 16385
<< pdiff >>
rect 7156 563 7275 722
rect 7156 517 7200 563
rect 7246 517 7275 563
rect 7156 359 7275 517
rect 7156 313 7200 359
rect 7246 313 7275 359
rect 7156 267 7275 313
rect 7395 267 7499 722
rect 7619 563 7723 722
rect 7619 517 7648 563
rect 7694 517 7723 563
rect 7619 359 7723 517
rect 7619 313 7648 359
rect 7694 313 7723 359
rect 7619 267 7723 313
rect 7843 267 7947 722
rect 8067 563 8185 722
rect 8067 517 8096 563
rect 8142 517 8185 563
rect 8067 359 8185 517
rect 8067 313 8096 359
rect 8142 313 8185 359
rect 8067 267 8185 313
<< pdiffc >>
rect 7200 517 7246 563
rect 7200 313 7246 359
rect 7648 517 7694 563
rect 7648 313 7694 359
rect 8096 517 8142 563
rect 8096 313 8142 359
<< psubdiff >>
rect 476 9109 18355 9169
rect 476 9063 882 9109
rect 928 9063 1040 9109
rect 1086 9063 1198 9109
rect 1244 9063 1356 9109
rect 1402 9063 1514 9109
rect 1560 9063 1672 9109
rect 1718 9063 1831 9109
rect 1877 9063 1989 9109
rect 2035 9063 2147 9109
rect 2193 9063 2305 9109
rect 2351 9063 2463 9109
rect 2509 9063 2621 9109
rect 2667 9063 2779 9109
rect 2825 9063 2937 9109
rect 2983 9063 3095 9109
rect 3141 9063 3254 9109
rect 3300 9063 3412 9109
rect 3458 9063 3570 9109
rect 3616 9063 3728 9109
rect 3774 9063 3886 9109
rect 3932 9063 4044 9109
rect 4090 9063 4202 9109
rect 4248 9063 4360 9109
rect 4406 9063 4518 9109
rect 4564 9063 4677 9109
rect 4723 9063 4835 9109
rect 4881 9063 4993 9109
rect 5039 9063 5151 9109
rect 5197 9063 5309 9109
rect 5355 9063 5467 9109
rect 5513 9063 5625 9109
rect 5671 9063 5783 9109
rect 5829 9063 5941 9109
rect 5987 9063 6100 9109
rect 6146 9063 6258 9109
rect 6304 9063 6416 9109
rect 6462 9063 6574 9109
rect 6620 9063 6732 9109
rect 6778 9063 6890 9109
rect 6936 9063 7048 9109
rect 7094 9063 7206 9109
rect 7252 9063 7364 9109
rect 7410 9063 7523 9109
rect 7569 9063 7681 9109
rect 7727 9063 7839 9109
rect 7885 9063 7997 9109
rect 8043 9063 8155 9109
rect 8201 9063 8313 9109
rect 8359 9063 8471 9109
rect 8517 9063 8629 9109
rect 8675 9063 8787 9109
rect 8833 9063 8946 9109
rect 8992 9063 9104 9109
rect 9150 9063 9262 9109
rect 9308 9063 9420 9109
rect 9466 9063 9578 9109
rect 9624 9063 9736 9109
rect 9782 9063 9894 9109
rect 9940 9063 10052 9109
rect 10098 9063 10210 9109
rect 10256 9063 10369 9109
rect 10415 9063 10527 9109
rect 10573 9063 10685 9109
rect 10731 9063 10843 9109
rect 10889 9063 11001 9109
rect 11047 9063 11159 9109
rect 11205 9063 11317 9109
rect 11363 9063 11475 9109
rect 11521 9063 11634 9109
rect 11680 9063 11792 9109
rect 11838 9063 11950 9109
rect 11996 9063 12108 9109
rect 12154 9063 12266 9109
rect 12312 9063 12424 9109
rect 12470 9063 12582 9109
rect 12628 9063 12740 9109
rect 12786 9063 12898 9109
rect 12944 9063 13057 9109
rect 13103 9063 13215 9109
rect 13261 9063 13373 9109
rect 13419 9063 13531 9109
rect 13577 9063 13689 9109
rect 13735 9063 13847 9109
rect 13893 9063 14005 9109
rect 14051 9063 14163 9109
rect 14209 9063 14321 9109
rect 14367 9063 14480 9109
rect 14526 9063 14638 9109
rect 14684 9063 14796 9109
rect 14842 9063 14954 9109
rect 15000 9063 15112 9109
rect 15158 9063 15270 9109
rect 15316 9063 15428 9109
rect 15474 9063 15586 9109
rect 15632 9063 15744 9109
rect 15790 9063 15903 9109
rect 15949 9063 16061 9109
rect 16107 9063 16219 9109
rect 16265 9063 16377 9109
rect 16423 9063 16535 9109
rect 16581 9063 16693 9109
rect 16739 9063 16851 9109
rect 16897 9063 17009 9109
rect 17055 9063 17167 9109
rect 17213 9063 17326 9109
rect 17372 9063 17484 9109
rect 17530 9063 17642 9109
rect 17688 9063 17800 9109
rect 17846 9063 17958 9109
rect 18004 9063 18116 9109
rect 18162 9063 18274 9109
rect 18320 9063 18355 9109
rect 476 9004 18355 9063
<< psubdiffcont >>
rect 882 9063 928 9109
rect 1040 9063 1086 9109
rect 1198 9063 1244 9109
rect 1356 9063 1402 9109
rect 1514 9063 1560 9109
rect 1672 9063 1718 9109
rect 1831 9063 1877 9109
rect 1989 9063 2035 9109
rect 2147 9063 2193 9109
rect 2305 9063 2351 9109
rect 2463 9063 2509 9109
rect 2621 9063 2667 9109
rect 2779 9063 2825 9109
rect 2937 9063 2983 9109
rect 3095 9063 3141 9109
rect 3254 9063 3300 9109
rect 3412 9063 3458 9109
rect 3570 9063 3616 9109
rect 3728 9063 3774 9109
rect 3886 9063 3932 9109
rect 4044 9063 4090 9109
rect 4202 9063 4248 9109
rect 4360 9063 4406 9109
rect 4518 9063 4564 9109
rect 4677 9063 4723 9109
rect 4835 9063 4881 9109
rect 4993 9063 5039 9109
rect 5151 9063 5197 9109
rect 5309 9063 5355 9109
rect 5467 9063 5513 9109
rect 5625 9063 5671 9109
rect 5783 9063 5829 9109
rect 5941 9063 5987 9109
rect 6100 9063 6146 9109
rect 6258 9063 6304 9109
rect 6416 9063 6462 9109
rect 6574 9063 6620 9109
rect 6732 9063 6778 9109
rect 6890 9063 6936 9109
rect 7048 9063 7094 9109
rect 7206 9063 7252 9109
rect 7364 9063 7410 9109
rect 7523 9063 7569 9109
rect 7681 9063 7727 9109
rect 7839 9063 7885 9109
rect 7997 9063 8043 9109
rect 8155 9063 8201 9109
rect 8313 9063 8359 9109
rect 8471 9063 8517 9109
rect 8629 9063 8675 9109
rect 8787 9063 8833 9109
rect 8946 9063 8992 9109
rect 9104 9063 9150 9109
rect 9262 9063 9308 9109
rect 9420 9063 9466 9109
rect 9578 9063 9624 9109
rect 9736 9063 9782 9109
rect 9894 9063 9940 9109
rect 10052 9063 10098 9109
rect 10210 9063 10256 9109
rect 10369 9063 10415 9109
rect 10527 9063 10573 9109
rect 10685 9063 10731 9109
rect 10843 9063 10889 9109
rect 11001 9063 11047 9109
rect 11159 9063 11205 9109
rect 11317 9063 11363 9109
rect 11475 9063 11521 9109
rect 11634 9063 11680 9109
rect 11792 9063 11838 9109
rect 11950 9063 11996 9109
rect 12108 9063 12154 9109
rect 12266 9063 12312 9109
rect 12424 9063 12470 9109
rect 12582 9063 12628 9109
rect 12740 9063 12786 9109
rect 12898 9063 12944 9109
rect 13057 9063 13103 9109
rect 13215 9063 13261 9109
rect 13373 9063 13419 9109
rect 13531 9063 13577 9109
rect 13689 9063 13735 9109
rect 13847 9063 13893 9109
rect 14005 9063 14051 9109
rect 14163 9063 14209 9109
rect 14321 9063 14367 9109
rect 14480 9063 14526 9109
rect 14638 9063 14684 9109
rect 14796 9063 14842 9109
rect 14954 9063 15000 9109
rect 15112 9063 15158 9109
rect 15270 9063 15316 9109
rect 15428 9063 15474 9109
rect 15586 9063 15632 9109
rect 15744 9063 15790 9109
rect 15903 9063 15949 9109
rect 16061 9063 16107 9109
rect 16219 9063 16265 9109
rect 16377 9063 16423 9109
rect 16535 9063 16581 9109
rect 16693 9063 16739 9109
rect 16851 9063 16897 9109
rect 17009 9063 17055 9109
rect 17167 9063 17213 9109
rect 17326 9063 17372 9109
rect 17484 9063 17530 9109
rect 17642 9063 17688 9109
rect 17800 9063 17846 9109
rect 17958 9063 18004 9109
rect 18116 9063 18162 9109
rect 18274 9063 18320 9109
<< polysilicon >>
rect 7429 1211 7566 1230
rect 7429 1071 7448 1211
rect 7494 1071 7566 1211
rect 7429 1052 7566 1071
rect 6352 758 6472 967
rect 7499 942 7566 1052
rect 7722 942 7842 971
rect 7174 872 7395 891
rect 7174 826 7193 872
rect 7239 826 7395 872
rect 7174 807 7395 826
rect 6246 683 6590 758
rect 7275 722 7395 807
rect 7499 876 7842 942
rect 7946 907 8066 971
rect 7946 891 8240 907
rect 7947 888 8240 891
rect 7499 820 7843 876
rect 7499 722 7619 820
rect 7723 722 7843 820
rect 7947 842 8081 888
rect 8221 842 8240 888
rect 7947 823 8240 842
rect 7947 722 8067 823
rect 6246 664 6366 683
rect 6470 664 6590 683
rect 6246 221 6366 240
rect 6470 221 6590 240
rect 6246 202 6590 221
rect 6246 156 6307 202
rect 6541 156 6590 202
rect 7275 194 7395 267
rect 7499 194 7619 267
rect 7723 194 7843 267
rect 7947 194 8067 267
rect 6246 137 6590 156
<< polycontact >>
rect 7448 1071 7494 1211
rect 7193 826 7239 872
rect 8081 842 8221 888
rect 6307 156 6541 202
<< metal1 >>
rect 392 16122 18614 16364
rect 399 9302 515 9303
rect 1071 9302 1187 9303
rect 1519 9302 1635 9303
rect 2191 9302 2307 9303
rect 2639 9302 2755 9303
rect 3311 9302 3427 9303
rect 3759 9302 3875 9303
rect 4431 9302 4547 9303
rect 4879 9302 4995 9303
rect 5551 9302 5667 9303
rect 5999 9302 6115 9303
rect 6671 9302 6787 9303
rect 7119 9302 7235 9303
rect 7791 9302 7907 9303
rect 8239 9302 8355 9303
rect 8911 9302 9027 9303
rect 9359 9302 9475 9303
rect 10031 9302 10147 9303
rect 10479 9302 10595 9303
rect 11151 9302 11267 9303
rect 11599 9302 11715 9303
rect 12271 9302 12387 9303
rect 12719 9302 12835 9303
rect 13391 9302 13507 9303
rect 13839 9302 13955 9303
rect 14511 9302 14627 9303
rect 14959 9302 15075 9303
rect 15630 9302 15747 9303
rect 16078 9302 16195 9303
rect 16750 9302 16867 9303
rect 17198 9302 17315 9303
rect 17870 9302 17987 9303
rect 18318 9302 18434 9303
rect 373 9109 18434 9302
rect 373 9063 882 9109
rect 928 9063 1040 9109
rect 1086 9063 1198 9109
rect 1244 9063 1356 9109
rect 1402 9063 1514 9109
rect 1560 9063 1672 9109
rect 1718 9063 1831 9109
rect 1877 9063 1989 9109
rect 2035 9063 2147 9109
rect 2193 9063 2305 9109
rect 2351 9063 2463 9109
rect 2509 9063 2621 9109
rect 2667 9063 2779 9109
rect 2825 9063 2937 9109
rect 2983 9063 3095 9109
rect 3141 9063 3254 9109
rect 3300 9063 3412 9109
rect 3458 9063 3570 9109
rect 3616 9063 3728 9109
rect 3774 9063 3886 9109
rect 3932 9063 4044 9109
rect 4090 9063 4202 9109
rect 4248 9063 4360 9109
rect 4406 9063 4518 9109
rect 4564 9063 4677 9109
rect 4723 9063 4835 9109
rect 4881 9063 4993 9109
rect 5039 9063 5151 9109
rect 5197 9063 5309 9109
rect 5355 9063 5467 9109
rect 5513 9063 5625 9109
rect 5671 9063 5783 9109
rect 5829 9063 5941 9109
rect 5987 9063 6100 9109
rect 6146 9063 6258 9109
rect 6304 9063 6416 9109
rect 6462 9063 6574 9109
rect 6620 9063 6732 9109
rect 6778 9063 6890 9109
rect 6936 9063 7048 9109
rect 7094 9063 7206 9109
rect 7252 9063 7364 9109
rect 7410 9063 7523 9109
rect 7569 9063 7681 9109
rect 7727 9063 7839 9109
rect 7885 9063 7997 9109
rect 8043 9063 8155 9109
rect 8201 9063 8313 9109
rect 8359 9063 8471 9109
rect 8517 9063 8629 9109
rect 8675 9063 8787 9109
rect 8833 9063 8946 9109
rect 8992 9063 9104 9109
rect 9150 9063 9262 9109
rect 9308 9063 9420 9109
rect 9466 9063 9578 9109
rect 9624 9063 9736 9109
rect 9782 9063 9894 9109
rect 9940 9063 10052 9109
rect 10098 9063 10210 9109
rect 10256 9063 10369 9109
rect 10415 9063 10527 9109
rect 10573 9063 10685 9109
rect 10731 9063 10843 9109
rect 10889 9063 11001 9109
rect 11047 9063 11159 9109
rect 11205 9063 11317 9109
rect 11363 9063 11475 9109
rect 11521 9063 11634 9109
rect 11680 9063 11792 9109
rect 11838 9063 11950 9109
rect 11996 9063 12108 9109
rect 12154 9063 12266 9109
rect 12312 9063 12424 9109
rect 12470 9063 12582 9109
rect 12628 9063 12740 9109
rect 12786 9063 12898 9109
rect 12944 9063 13057 9109
rect 13103 9063 13215 9109
rect 13261 9063 13373 9109
rect 13419 9063 13531 9109
rect 13577 9063 13689 9109
rect 13735 9063 13847 9109
rect 13893 9063 14005 9109
rect 14051 9063 14163 9109
rect 14209 9063 14321 9109
rect 14367 9063 14480 9109
rect 14526 9063 14638 9109
rect 14684 9063 14796 9109
rect 14842 9063 14954 9109
rect 15000 9063 15112 9109
rect 15158 9063 15270 9109
rect 15316 9063 15428 9109
rect 15474 9063 15586 9109
rect 15632 9063 15744 9109
rect 15790 9063 15903 9109
rect 15949 9063 16061 9109
rect 16107 9063 16219 9109
rect 16265 9063 16377 9109
rect 16423 9063 16535 9109
rect 16581 9063 16693 9109
rect 16739 9063 16851 9109
rect 16897 9063 17009 9109
rect 17055 9063 17167 9109
rect 17213 9063 17326 9109
rect 17372 9063 17484 9109
rect 17530 9063 17642 9109
rect 17688 9063 17800 9109
rect 17846 9063 17958 9109
rect 18004 9063 18116 9109
rect 18162 9063 18274 9109
rect 18320 9063 18434 9109
rect 373 8697 18434 9063
rect 1242 4508 1371 5054
rect 2933 4379 3062 4420
rect 2933 4327 2972 4379
rect 3024 4327 3062 4379
rect 2933 4286 3062 4327
rect 4623 4177 4752 4218
rect 4623 4125 4662 4177
rect 4714 4125 4752 4177
rect 4623 4084 4752 4125
rect 1755 3975 1884 4016
rect 1755 3923 1794 3975
rect 1846 3923 1884 3975
rect 1755 3882 1884 3923
rect 3446 3773 3575 3814
rect 3446 3721 3485 3773
rect 3537 3721 3575 3773
rect 3446 3680 3575 3721
rect 5137 3572 5266 3613
rect 5137 3520 5176 3572
rect 5228 3520 5266 3572
rect 5137 3479 5266 3520
rect 5399 196 5528 2118
rect 6242 1618 6358 1690
rect 6243 1357 6358 1618
rect 6242 1356 6358 1357
rect 7404 1366 7528 1406
rect 6241 1316 6365 1356
rect 6241 1264 6277 1316
rect 6329 1264 6365 1316
rect 6241 1098 6365 1264
rect 7404 1314 7440 1366
rect 7492 1314 7528 1366
rect 7404 1211 7528 1314
rect 6241 1046 6277 1098
rect 6329 1046 6365 1098
rect 6241 1006 6365 1046
rect 5621 874 5745 907
rect 6467 874 6582 1180
rect 7404 1148 7448 1211
rect 7404 1096 7440 1148
rect 7404 1071 7448 1096
rect 7494 1071 7528 1211
rect 7404 1056 7528 1071
rect 7647 1010 7693 1717
rect 7871 915 7917 1316
rect 8095 1128 12303 1724
rect 8095 1010 8141 1128
rect 5619 867 6582 874
rect 5619 815 5657 867
rect 5709 815 6582 867
rect 7069 891 7353 903
rect 7069 839 7081 891
rect 7341 839 7353 891
rect 7069 827 7193 839
rect 7182 826 7193 827
rect 7239 827 7353 839
rect 7239 826 7250 827
rect 7182 815 7250 826
rect 5619 740 6582 815
rect 7631 795 7917 915
rect 8040 891 8324 903
rect 8040 839 8052 891
rect 8312 839 8324 891
rect 8040 827 8324 839
rect 5621 649 5745 740
rect 5621 597 5657 649
rect 5709 597 5745 649
rect 5621 557 5745 597
rect 5850 623 5974 640
rect 5850 600 6217 623
rect 5850 548 5886 600
rect 5938 548 6217 600
rect 5850 382 6217 548
rect 5850 330 5886 382
rect 5938 330 6217 382
rect 6395 378 6441 740
rect 6877 623 7001 658
rect 6619 618 7281 623
rect 6619 566 6913 618
rect 6965 566 7281 618
rect 6619 563 7281 566
rect 6619 517 7200 563
rect 7246 517 7281 563
rect 6619 400 7281 517
rect 5850 281 6217 330
rect 6619 348 6913 400
rect 6965 359 7281 400
rect 6965 348 7200 359
rect 6619 313 7200 348
rect 7246 313 7281 359
rect 6619 281 7281 313
rect 7165 276 7281 281
rect 7631 563 7710 795
rect 7631 517 7648 563
rect 7694 517 7710 563
rect 7631 359 7710 517
rect 7631 313 7648 359
rect 7694 313 7710 359
rect 6296 202 6552 213
rect 6296 196 6307 202
rect 5399 156 6307 196
rect 6541 196 6552 202
rect 7631 196 7710 313
rect 8061 563 12088 681
rect 8061 517 8096 563
rect 8142 517 12088 563
rect 8061 359 12088 517
rect 8061 313 8096 359
rect 8142 313 12088 359
rect 8061 276 12088 313
rect 6541 156 7710 196
rect 5399 76 7710 156
<< via1 >>
rect 2972 4327 3024 4379
rect 4662 4125 4714 4177
rect 1794 3923 1846 3975
rect 3485 3721 3537 3773
rect 5176 3520 5228 3572
rect 6277 1264 6329 1316
rect 7440 1314 7492 1366
rect 6277 1046 6329 1098
rect 7440 1096 7448 1148
rect 7448 1096 7492 1148
rect 5657 815 5709 867
rect 7081 872 7341 891
rect 7081 839 7193 872
rect 7193 839 7239 872
rect 7239 839 7341 872
rect 8052 888 8312 891
rect 8052 842 8081 888
rect 8081 842 8221 888
rect 8221 842 8312 888
rect 8052 839 8312 842
rect 5657 597 5709 649
rect 5886 548 5938 600
rect 5886 330 5938 382
rect 6913 566 6965 618
rect 6913 348 6965 400
<< metal2 >>
rect 8679 14374 8808 14413
rect 8679 14318 8716 14374
rect 8772 14318 8808 14374
rect 8679 14279 8808 14318
rect 9127 14374 9256 14413
rect 9127 14318 9164 14374
rect 9220 14318 9256 14374
rect 9127 14279 9256 14318
rect 17640 14374 17769 14413
rect 17640 14318 17676 14374
rect 17732 14318 17769 14374
rect 17640 14279 17769 14318
rect 18088 14374 18217 14413
rect 18088 14318 18124 14374
rect 18180 14318 18217 14374
rect 18088 14279 18217 14318
rect 7560 14034 7689 14073
rect 7560 13978 7597 14034
rect 7653 13978 7689 14034
rect 7560 13939 7689 13978
rect 8007 14034 8136 14073
rect 8007 13978 8044 14034
rect 8100 13978 8136 14034
rect 8007 13939 8136 13978
rect 16520 14034 16649 14073
rect 16520 13978 16556 14034
rect 16612 13978 16649 14034
rect 16520 13939 16649 13978
rect 16968 14034 17097 14073
rect 16968 13978 17004 14034
rect 17060 13978 17097 14034
rect 16968 13939 17097 13978
rect 6440 13693 6569 13732
rect 6440 13637 6477 13693
rect 6533 13637 6569 13693
rect 6440 13598 6569 13637
rect 6888 13693 7017 13732
rect 6888 13637 6925 13693
rect 6981 13637 7017 13693
rect 6888 13598 7017 13637
rect 15400 13693 15529 13732
rect 15400 13637 15436 13693
rect 15492 13637 15529 13693
rect 15400 13598 15529 13637
rect 15848 13693 15977 13732
rect 15848 13637 15884 13693
rect 15940 13637 15977 13693
rect 15848 13598 15977 13637
rect 5320 13353 5449 13392
rect 5320 13297 5357 13353
rect 5413 13297 5449 13353
rect 5320 13258 5449 13297
rect 5768 13353 5897 13392
rect 5768 13297 5805 13353
rect 5861 13297 5897 13353
rect 5768 13258 5897 13297
rect 14280 13353 14409 13392
rect 14280 13297 14316 13353
rect 14372 13297 14409 13353
rect 14280 13258 14409 13297
rect 14728 13353 14857 13392
rect 14728 13297 14764 13353
rect 14820 13297 14857 13353
rect 14728 13258 14857 13297
rect 4200 13013 4329 13052
rect 4200 12957 4237 13013
rect 4293 12957 4329 13013
rect 4200 12918 4329 12957
rect 4648 13013 4777 13052
rect 4648 12957 4685 13013
rect 4741 12957 4777 13013
rect 4648 12918 4777 12957
rect 13160 13013 13289 13052
rect 13160 12957 13196 13013
rect 13252 12957 13289 13013
rect 13160 12918 13289 12957
rect 13608 13013 13737 13052
rect 13608 12957 13644 13013
rect 13700 12957 13737 13013
rect 13608 12918 13737 12957
rect 3080 12673 3209 12712
rect 3080 12617 3117 12673
rect 3173 12617 3209 12673
rect 3080 12578 3209 12617
rect 3528 12673 3657 12712
rect 3528 12617 3565 12673
rect 3621 12617 3657 12673
rect 3528 12578 3657 12617
rect 12040 12673 12169 12712
rect 12040 12617 12076 12673
rect 12132 12617 12169 12673
rect 12040 12578 12169 12617
rect 12488 12673 12617 12712
rect 12488 12617 12524 12673
rect 12580 12617 12617 12673
rect 12488 12578 12617 12617
rect 1960 12333 2089 12372
rect 1960 12277 1997 12333
rect 2053 12277 2089 12333
rect 1960 12238 2089 12277
rect 2408 12333 2537 12372
rect 2408 12277 2445 12333
rect 2501 12277 2537 12333
rect 2408 12238 2537 12277
rect 10920 12333 11049 12372
rect 10920 12277 10956 12333
rect 11012 12277 11049 12333
rect 10920 12238 11049 12277
rect 11368 12333 11497 12372
rect 11368 12277 11404 12333
rect 11460 12277 11497 12333
rect 11368 12238 11497 12277
rect 840 11993 969 12032
rect 840 11937 877 11993
rect 933 11937 969 11993
rect 840 11898 969 11937
rect 1288 11993 1417 12032
rect 1288 11937 1325 11993
rect 1381 11937 1417 11993
rect 1288 11898 1417 11937
rect 9800 11993 9929 12032
rect 9800 11937 9836 11993
rect 9892 11937 9929 11993
rect 9800 11898 9929 11937
rect 10248 11993 10377 12032
rect 10248 11937 10284 11993
rect 10340 11937 10377 11993
rect 10248 11898 10377 11937
rect 409 11592 534 11631
rect 409 11536 444 11592
rect 500 11536 534 11592
rect 11145 11608 11270 11647
rect 11145 11552 11180 11608
rect 11236 11552 11270 11608
rect 11145 11538 11270 11552
rect 409 11374 534 11536
rect 9367 11499 9707 11538
rect 9367 11443 9403 11499
rect 9459 11443 9615 11499
rect 9671 11443 9707 11499
rect 409 11318 444 11374
rect 500 11318 534 11374
rect 409 11280 534 11318
rect 1528 11290 1868 11329
rect 1528 11234 1564 11290
rect 1620 11234 1776 11290
rect 1832 11234 1868 11290
rect 1528 11195 1868 11234
rect 2648 11062 2777 11413
rect 2648 11008 2684 11062
rect 2649 11006 2684 11008
rect 2740 11008 2777 11062
rect 2740 11006 2774 11008
rect 2649 10844 2774 11006
rect 3768 10912 3897 11413
rect 2649 10788 2684 10844
rect 2740 10788 2774 10844
rect 2649 10750 2774 10788
rect 3767 10873 4107 10912
rect 3767 10817 3803 10873
rect 3859 10817 4015 10873
rect 4071 10817 4107 10873
rect 3767 10778 4107 10817
rect 4888 10704 5017 11413
rect 4782 10665 5122 10704
rect 4782 10609 4818 10665
rect 4874 10609 5030 10665
rect 5086 10609 5122 10665
rect 4782 10570 5122 10609
rect 6008 10495 6137 11413
rect 5902 10456 6242 10495
rect 5902 10400 5938 10456
rect 5994 10400 6150 10456
rect 6206 10400 6242 10456
rect 5902 10361 6242 10400
rect 7128 10287 7257 11413
rect 7720 10456 8060 10495
rect 7720 10400 7756 10456
rect 7812 10400 7968 10456
rect 8024 10400 8060 10456
rect 7720 10361 8060 10400
rect 6829 10286 7257 10287
rect 6741 10248 7257 10286
rect 6741 10192 6865 10248
rect 6921 10192 7077 10248
rect 7133 10192 7257 10248
rect 6741 10153 7257 10192
rect 6192 10039 6532 10078
rect 6192 9983 6228 10039
rect 6284 9983 6440 10039
rect 6496 9983 6532 10039
rect 6192 9944 6532 9983
rect 6297 8727 6426 9944
rect 6741 8727 6870 10153
rect 7931 8727 8060 10361
rect 8248 10078 8377 11413
rect 9367 11404 9707 11443
rect 11144 11390 11273 11538
rect 11144 11334 11180 11390
rect 11236 11334 11273 11390
rect 10487 11290 10827 11329
rect 10487 11234 10523 11290
rect 10579 11234 10735 11290
rect 10791 11234 10827 11290
rect 10487 11195 10827 11234
rect 10021 11100 10150 11121
rect 10021 11082 10151 11100
rect 10021 11026 10058 11082
rect 10114 11026 10151 11082
rect 10021 10987 10151 11026
rect 9354 10873 9694 10912
rect 9354 10817 9390 10873
rect 9446 10817 9602 10873
rect 9658 10817 9694 10873
rect 9354 10778 9694 10817
rect 8671 10665 9011 10704
rect 8671 10609 8707 10665
rect 8763 10609 8919 10665
rect 8975 10609 9011 10665
rect 8671 10570 9011 10609
rect 8247 10039 8587 10078
rect 8247 9983 8283 10039
rect 8339 9983 8495 10039
rect 8551 9983 8587 10039
rect 8247 9944 8587 9983
rect 8777 9640 8906 10570
rect 8375 9507 8906 9640
rect 8375 8727 8504 9507
rect 9565 8727 9694 10778
rect 10022 9516 10151 10987
rect 10009 9382 10151 9516
rect 10487 9541 10616 11195
rect 11144 9905 11273 11334
rect 11607 11128 11736 11413
rect 11607 11127 11737 11128
rect 11607 11089 11946 11127
rect 11607 11033 11643 11089
rect 11699 11033 11855 11089
rect 11911 11033 11946 11089
rect 11607 10994 11946 11033
rect 12727 11112 12856 11413
rect 12727 11056 12764 11112
rect 12820 11056 12856 11112
rect 12727 10894 12856 11056
rect 12727 10838 12764 10894
rect 12820 10838 12856 10894
rect 12727 10799 12856 10838
rect 13847 10903 13976 11413
rect 13847 10847 13884 10903
rect 13940 10847 13976 10903
rect 13847 10685 13976 10847
rect 13847 10629 13884 10685
rect 13940 10629 13976 10685
rect 13847 10590 13976 10629
rect 14967 10694 15096 11413
rect 14967 10638 15004 10694
rect 15060 10638 15096 10694
rect 14967 10476 15096 10638
rect 14967 10420 15004 10476
rect 15060 10420 15096 10476
rect 14967 10382 15096 10420
rect 16087 10486 16216 11413
rect 16087 10430 16124 10486
rect 16180 10430 16216 10486
rect 16087 10268 16216 10430
rect 16087 10212 16124 10268
rect 16180 10212 16216 10268
rect 16087 10173 16216 10212
rect 17207 10277 17336 11631
rect 17207 10221 17244 10277
rect 17300 10221 17336 10277
rect 17207 10059 17336 10221
rect 17207 10003 17244 10059
rect 17300 10003 17336 10059
rect 17207 9965 17336 10003
rect 11144 9772 11772 9905
rect 10487 9540 10617 9541
rect 10487 9407 11328 9540
rect 10009 8727 10138 9382
rect 11199 8727 11328 9407
rect 11643 8727 11772 9772
rect 1756 4016 1885 5054
rect 2933 4379 3062 5054
rect 2933 4327 2972 4379
rect 3024 4327 3062 4379
rect 2933 4286 3062 4327
rect 1755 3975 1885 4016
rect 1755 3923 1794 3975
rect 1846 3923 1885 3975
rect 1755 3903 1885 3923
rect 1755 3882 1884 3903
rect 3447 3814 3576 5054
rect 4624 4218 4753 5054
rect 4623 4177 4753 4218
rect 4623 4125 4662 4177
rect 4714 4125 4753 4177
rect 4623 4105 4753 4125
rect 4623 4084 4752 4105
rect 3446 3773 3576 3814
rect 3446 3721 3485 3773
rect 3537 3721 3576 3773
rect 3446 3701 3576 3721
rect 3446 3680 3575 3701
rect 5138 3613 5267 4823
rect 5137 3572 5267 3613
rect 5137 3520 5176 3572
rect 5228 3520 5267 3572
rect 5137 3499 5267 3520
rect 5137 3479 5266 3499
rect 5399 2642 5748 2776
rect 5619 867 5748 2642
rect 7402 1366 7531 1406
rect 6241 1318 6366 1357
rect 6241 1262 6275 1318
rect 6331 1262 6366 1318
rect 7402 1314 7440 1366
rect 7492 1314 7531 1366
rect 7402 1273 7531 1314
rect 6241 1100 6366 1262
rect 6241 1044 6275 1100
rect 6331 1044 6366 1100
rect 7404 1148 7528 1273
rect 7404 1096 7440 1148
rect 7492 1096 7528 1148
rect 7404 1056 7528 1096
rect 6241 1006 6366 1044
rect 5619 815 5657 867
rect 5709 815 5748 867
rect 7069 891 8324 903
rect 7069 839 7081 891
rect 7341 839 8052 891
rect 8312 839 8324 891
rect 7069 827 8324 839
rect 1811 607 1940 740
rect 3502 607 3631 740
rect 5193 607 5322 740
rect 5619 649 5748 815
rect 5619 597 5657 649
rect 5709 597 5748 649
rect 5619 557 5748 597
rect 5850 602 5975 641
rect 5850 546 5884 602
rect 5940 546 5975 602
rect 5850 384 5975 546
rect 5850 328 5884 384
rect 5940 328 5975 384
rect 5850 290 5975 328
rect 6877 620 7002 659
rect 6877 564 6911 620
rect 6967 564 7002 620
rect 6877 402 7002 564
rect 6877 346 6911 402
rect 6967 346 7002 402
rect 6877 308 7002 346
<< via2 >>
rect 8716 14318 8772 14374
rect 9164 14318 9220 14374
rect 17676 14318 17732 14374
rect 18124 14318 18180 14374
rect 7597 13978 7653 14034
rect 8044 13978 8100 14034
rect 16556 13978 16612 14034
rect 17004 13978 17060 14034
rect 6477 13637 6533 13693
rect 6925 13637 6981 13693
rect 15436 13637 15492 13693
rect 15884 13637 15940 13693
rect 5357 13297 5413 13353
rect 5805 13297 5861 13353
rect 14316 13297 14372 13353
rect 14764 13297 14820 13353
rect 4237 12957 4293 13013
rect 4685 12957 4741 13013
rect 13196 12957 13252 13013
rect 13644 12957 13700 13013
rect 3117 12617 3173 12673
rect 3565 12617 3621 12673
rect 12076 12617 12132 12673
rect 12524 12617 12580 12673
rect 1997 12277 2053 12333
rect 2445 12277 2501 12333
rect 10956 12277 11012 12333
rect 11404 12277 11460 12333
rect 877 11937 933 11993
rect 1325 11937 1381 11993
rect 9836 11937 9892 11993
rect 10284 11937 10340 11993
rect 444 11536 500 11592
rect 11180 11552 11236 11608
rect 9403 11443 9459 11499
rect 9615 11443 9671 11499
rect 444 11318 500 11374
rect 1564 11234 1620 11290
rect 1776 11234 1832 11290
rect 2684 11006 2740 11062
rect 2684 10788 2740 10844
rect 3803 10817 3859 10873
rect 4015 10817 4071 10873
rect 4818 10609 4874 10665
rect 5030 10609 5086 10665
rect 5938 10400 5994 10456
rect 6150 10400 6206 10456
rect 7756 10400 7812 10456
rect 7968 10400 8024 10456
rect 6865 10192 6921 10248
rect 7077 10192 7133 10248
rect 6228 9983 6284 10039
rect 6440 9983 6496 10039
rect 11180 11334 11236 11390
rect 10523 11234 10579 11290
rect 10735 11234 10791 11290
rect 10058 11026 10114 11082
rect 9390 10817 9446 10873
rect 9602 10817 9658 10873
rect 8707 10609 8763 10665
rect 8919 10609 8975 10665
rect 8283 9983 8339 10039
rect 8495 9983 8551 10039
rect 11643 11033 11699 11089
rect 11855 11033 11911 11089
rect 12764 11056 12820 11112
rect 12764 10838 12820 10894
rect 13884 10847 13940 10903
rect 13884 10629 13940 10685
rect 15004 10638 15060 10694
rect 15004 10420 15060 10476
rect 16124 10430 16180 10486
rect 16124 10212 16180 10268
rect 17244 10221 17300 10277
rect 17244 10003 17300 10059
rect 6275 1316 6331 1318
rect 6275 1264 6277 1316
rect 6277 1264 6329 1316
rect 6329 1264 6331 1316
rect 6275 1262 6331 1264
rect 6275 1098 6331 1100
rect 6275 1046 6277 1098
rect 6277 1046 6329 1098
rect 6329 1046 6331 1098
rect 6275 1044 6331 1046
rect 5884 600 5940 602
rect 5884 548 5886 600
rect 5886 548 5938 600
rect 5938 548 5940 600
rect 5884 546 5940 548
rect 5884 382 5940 384
rect 5884 330 5886 382
rect 5886 330 5938 382
rect 5938 330 5940 382
rect 5884 328 5940 330
rect 6911 618 6967 620
rect 6911 566 6913 618
rect 6913 566 6965 618
rect 6965 566 6967 618
rect 6911 564 6967 566
rect 6911 400 6967 402
rect 6911 348 6913 400
rect 6913 348 6965 400
rect 6965 348 6967 400
rect 6911 346 6967 348
<< metal3 >>
rect 179 14374 9257 14460
rect 17640 14413 26678 14460
rect 179 14318 8716 14374
rect 8772 14318 9164 14374
rect 9220 14318 9257 14374
rect 179 14231 9257 14318
rect 17639 14374 26678 14413
rect 17639 14318 17676 14374
rect 17732 14318 18124 14374
rect 18180 14318 26678 14374
rect 17639 14279 26678 14318
rect 17640 14231 26678 14279
rect 179 14034 8139 14120
rect 16520 14073 26678 14120
rect 179 13978 7597 14034
rect 7653 13978 8044 14034
rect 8100 13978 8139 14034
rect 179 13891 8139 13978
rect 16519 14034 26678 14073
rect 16519 13978 16556 14034
rect 16612 13978 17004 14034
rect 17060 13978 26678 14034
rect 16519 13939 26678 13978
rect 16520 13891 26678 13939
rect 179 13732 7017 13780
rect 15400 13732 26678 13780
rect 179 13693 7018 13732
rect 179 13637 6477 13693
rect 6533 13637 6925 13693
rect 6981 13637 7018 13693
rect 179 13598 7018 13637
rect 15399 13693 26678 13732
rect 15399 13637 15436 13693
rect 15492 13637 15884 13693
rect 15940 13637 26678 13693
rect 15399 13598 26678 13637
rect 179 13551 7017 13598
rect 15400 13551 26678 13598
rect 179 13392 5897 13440
rect 14280 13392 26678 13440
rect 179 13353 5898 13392
rect 179 13297 5357 13353
rect 5413 13297 5805 13353
rect 5861 13297 5898 13353
rect 179 13258 5898 13297
rect 14279 13353 26678 13392
rect 14279 13297 14316 13353
rect 14372 13297 14764 13353
rect 14820 13297 26678 13353
rect 14279 13258 26678 13297
rect 179 13211 5897 13258
rect 14280 13211 26678 13258
rect 179 13052 4777 13100
rect 13160 13052 26678 13100
rect 179 13013 4778 13052
rect 179 12957 4237 13013
rect 4293 12957 4685 13013
rect 4741 12957 4778 13013
rect 179 12918 4778 12957
rect 13159 13013 26678 13052
rect 13159 12957 13196 13013
rect 13252 12957 13644 13013
rect 13700 12957 26678 13013
rect 13159 12918 26678 12957
rect 179 12871 4777 12918
rect 13160 12871 26678 12918
rect 179 12712 3657 12760
rect 12040 12712 26678 12760
rect 179 12673 3658 12712
rect 179 12617 3117 12673
rect 3173 12617 3565 12673
rect 3621 12617 3658 12673
rect 179 12578 3658 12617
rect 12039 12673 26678 12712
rect 12039 12617 12076 12673
rect 12132 12617 12524 12673
rect 12580 12617 26678 12673
rect 12039 12578 26678 12617
rect 179 12531 3657 12578
rect 12040 12531 26678 12578
rect 179 12372 2537 12420
rect 179 12333 2538 12372
rect 179 12277 1997 12333
rect 2053 12277 2445 12333
rect 2501 12277 2538 12333
rect 179 12238 2538 12277
rect 10918 12333 26678 12420
rect 10918 12277 10956 12333
rect 11012 12277 11404 12333
rect 11460 12277 26678 12333
rect 179 12191 2537 12238
rect 10918 12191 26678 12277
rect 179 12032 1417 12080
rect 9800 12032 26678 12080
rect 179 11993 1418 12032
rect 179 11937 877 11993
rect 933 11937 1325 11993
rect 1381 11937 1418 11993
rect 179 11898 1418 11937
rect 9799 11993 26678 12032
rect 9799 11937 9836 11993
rect 9892 11937 10284 11993
rect 10340 11937 26678 11993
rect 9799 11898 26678 11937
rect 179 11851 1417 11898
rect 9800 11851 26678 11898
rect 409 11592 535 11631
rect 409 11536 444 11592
rect 500 11536 535 11592
rect 11145 11608 11271 11647
rect 11145 11552 11180 11608
rect 11236 11552 11271 11608
rect 409 11517 535 11536
rect 9367 11517 9707 11538
rect 11145 11517 11271 11552
rect 409 11499 11273 11517
rect 409 11443 9403 11499
rect 9459 11443 9615 11499
rect 9671 11443 11273 11499
rect 409 11425 11273 11443
rect 409 11374 535 11425
rect 9367 11404 9707 11425
rect 409 11318 444 11374
rect 500 11318 535 11374
rect 11145 11390 11271 11425
rect 11145 11334 11180 11390
rect 11236 11334 11271 11390
rect 409 11279 535 11318
rect 1528 11309 1868 11329
rect 10487 11309 10827 11329
rect 1528 11290 10827 11309
rect 11145 11295 11271 11334
rect 1528 11234 1564 11290
rect 1620 11234 1776 11290
rect 1832 11234 10523 11290
rect 10579 11234 10735 11290
rect 10791 11234 10827 11290
rect 1528 11216 10827 11234
rect 1528 11195 1868 11216
rect 10487 11195 10827 11216
rect 2649 11100 2775 11101
rect 10021 11100 10151 11121
rect 11607 11100 11947 11127
rect 2648 11089 11947 11100
rect 2648 11082 11643 11089
rect 2648 11062 10058 11082
rect 2648 11008 2684 11062
rect 2649 11006 2684 11008
rect 2740 11026 10058 11062
rect 10114 11033 11643 11082
rect 11699 11033 11855 11089
rect 11911 11033 11947 11089
rect 10114 11026 11947 11033
rect 2740 11008 11947 11026
rect 2740 11006 2775 11008
rect 2649 10844 2775 11006
rect 10021 10987 10151 11008
rect 11607 10994 11947 11008
rect 12729 11112 12855 11151
rect 12729 11056 12764 11112
rect 12820 11056 12855 11112
rect 2649 10788 2684 10844
rect 2740 10788 2775 10844
rect 2649 10749 2775 10788
rect 3767 10892 4107 10912
rect 9354 10892 9694 10912
rect 12729 10894 12855 11056
rect 12729 10892 12764 10894
rect 3767 10873 12764 10892
rect 3767 10817 3803 10873
rect 3859 10817 4015 10873
rect 4071 10817 9390 10873
rect 9446 10817 9602 10873
rect 9658 10838 12764 10873
rect 12820 10892 12855 10894
rect 13849 10903 13975 10942
rect 12820 10838 12856 10892
rect 9658 10817 12856 10838
rect 3767 10799 12856 10817
rect 13849 10847 13884 10903
rect 13940 10847 13975 10903
rect 3767 10778 4107 10799
rect 9354 10778 9694 10799
rect 4782 10683 5122 10704
rect 8671 10683 9011 10704
rect 13849 10685 13975 10847
rect 13849 10683 13884 10685
rect 4782 10665 13884 10683
rect 4782 10609 4818 10665
rect 4874 10609 5030 10665
rect 5086 10609 8707 10665
rect 8763 10609 8919 10665
rect 8975 10629 13884 10665
rect 13940 10683 13975 10685
rect 14969 10694 15095 10733
rect 13940 10629 13976 10683
rect 8975 10609 13976 10629
rect 4782 10590 13976 10609
rect 14969 10638 15004 10694
rect 15060 10638 15095 10694
rect 4782 10570 5122 10590
rect 8671 10570 9011 10590
rect 5902 10475 6242 10495
rect 7720 10475 8060 10495
rect 14969 10476 15095 10638
rect 14969 10475 15004 10476
rect 5902 10456 15004 10475
rect 5902 10400 5938 10456
rect 5994 10400 6150 10456
rect 6206 10400 7756 10456
rect 7812 10400 7968 10456
rect 8024 10420 15004 10456
rect 15060 10475 15095 10476
rect 16089 10486 16215 10525
rect 15060 10420 15096 10475
rect 8024 10400 15096 10420
rect 5902 10382 15096 10400
rect 16089 10430 16124 10486
rect 16180 10430 16215 10486
rect 5902 10361 6242 10382
rect 7720 10361 8060 10382
rect 14969 10381 15095 10382
rect 6829 10266 7169 10287
rect 16089 10268 16215 10430
rect 16089 10266 16124 10268
rect 6829 10248 16124 10266
rect 6829 10192 6865 10248
rect 6921 10192 7077 10248
rect 7133 10212 16124 10248
rect 16180 10266 16215 10268
rect 17209 10277 17335 10316
rect 16180 10212 16216 10266
rect 7133 10192 16216 10212
rect 6829 10173 16216 10192
rect 17209 10221 17244 10277
rect 17300 10221 17335 10277
rect 6829 10153 7169 10173
rect 6192 10057 6532 10078
rect 8247 10057 8587 10078
rect 17209 10059 17335 10221
rect 17209 10057 17244 10059
rect 6192 10039 17244 10057
rect 6192 9983 6228 10039
rect 6284 9983 6440 10039
rect 6496 9983 8283 10039
rect 8339 9983 8495 10039
rect 8551 10003 17244 10039
rect 17300 10057 17335 10059
rect 17300 10003 17336 10057
rect 8551 9983 17336 10003
rect 6192 9965 17336 9983
rect 6192 9944 6532 9965
rect 8247 9944 8587 9965
rect 17209 9964 17335 9965
rect 384 7972 12446 9232
rect 419 2629 5869 3311
rect 443 1473 5471 2381
rect 5766 1318 12303 1733
rect 5766 1302 6275 1318
rect 4777 1262 6275 1302
rect 6331 1262 12303 1318
rect 4777 1100 12303 1262
rect 4777 1044 6275 1100
rect 6331 1044 12303 1100
rect 4777 906 12303 1044
rect 5694 620 12299 675
rect 5694 602 6911 620
rect 5694 546 5884 602
rect 5940 564 6911 602
rect 6967 564 12299 620
rect 5940 546 12299 564
rect 5694 402 12299 546
rect 5694 384 6911 402
rect 5694 328 5884 384
rect 5940 346 6911 384
rect 6967 346 12299 402
rect 5940 328 12299 346
rect 5694 226 12299 328
use M1_NWELL$$47634476_256x8m81  M1_NWELL$$47634476_256x8m81_0
timestamp 1666464484
transform 1 0 9487 0 1 16304
box -9233 -228 9233 228
use M1_NWELL$$47635500_256x8m81  M1_NWELL$$47635500_256x8m81_0
timestamp 1666464484
transform 1 0 10211 0 1 442
box -2039 -309 2039 309
use M1_POLY24310590878126_256x8m81  M1_POLY24310590878126_256x8m81_0
timestamp 1666464484
transform 1 0 6424 0 1 179
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1666464484
transform 1 0 7216 0 1 849
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1666464484
transform 0 -1 8151 1 0 865
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_1
timestamp 1666464484
transform 1 0 7471 0 1 1141
box 0 0 1 1
use M1_PSUB$$47114284_256x8m81  M1_PSUB$$47114284_256x8m81_0
timestamp 1666464484
transform 1 0 10240 0 1 1283
box -1898 -164 1898 164
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1666464484
transform -1 0 7466 0 1 1231
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1666464484
transform -1 0 5683 0 1 732
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1666464484
transform -1 0 6303 0 1 1181
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1666464484
transform -1 0 6939 0 1 483
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1666464484
transform -1 0 5912 0 1 465
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_0
timestamp 1666464484
transform -1 0 5202 0 1 3546
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_1
timestamp 1666464484
transform -1 0 4688 0 1 4151
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_2
timestamp 1666464484
transform -1 0 1820 0 1 3949
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_3
timestamp 1666464484
transform -1 0 3511 0 1 3747
box 0 0 1 1
use M2_M1$$46894124_256x8m81  M2_M1$$46894124_256x8m81_4
timestamp 1666464484
transform -1 0 2998 0 1 4353
box 0 0 1 1
use M2_M1$$47630380_256x8m81  M2_M1$$47630380_256x8m81_0
timestamp 1666464484
transform -1 0 10023 0 1 478
box -1962 -176 1962 176
use M2_M1$$47631404_256x8m81  M2_M1$$47631404_256x8m81_0
timestamp 1666464484
transform -1 0 10157 0 1 1313
box -1857 -176 1857 176
use M2_M14310590878145_256x8m81  M2_M14310590878145_256x8m81_0
timestamp 1666464484
transform 1 0 7211 0 1 865
box 0 0 1 1
use M2_M14310590878145_256x8m81  M2_M14310590878145_256x8m81_1
timestamp 1666464484
transform 1 0 8182 0 1 865
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_0
timestamp 1666464484
transform -1 0 6303 0 1 1181
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_1
timestamp 1666464484
transform -1 0 6939 0 1 483
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_2
timestamp 1666464484
transform -1 0 5912 0 1 465
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_3
timestamp 1666464484
transform 1 0 2712 0 1 10925
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_4
timestamp 1666464484
transform 1 0 472 0 1 11455
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_5
timestamp 1666464484
transform 1 0 11208 0 1 11471
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_6
timestamp 1666464484
transform 1 0 12792 0 1 10975
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_7
timestamp 1666464484
transform 1 0 13912 0 1 10766
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_8
timestamp 1666464484
transform 1 0 15032 0 1 10557
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_9
timestamp 1666464484
transform 1 0 16152 0 1 10349
box 0 0 1 1
use M3_M2$$43368492_256x8m81_0  M3_M2$$43368492_256x8m81_0_10
timestamp 1666464484
transform 1 0 17272 0 1 10140
box 0 0 1 1
use M3_M2$$43368492_R90_256x8m81  M3_M2$$43368492_R90_256x8m81_0
timestamp 1666464484
transform 0 -1 10657 1 0 11262
box 0 0 1 1
use M3_M2$$43368492_R270_256x8m81  M3_M2$$43368492_R270_256x8m81_0
timestamp 1666464484
transform 0 1 11777 -1 0 11061
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_0
timestamp 1666464484
transform 1 0 8841 0 1 10637
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_1
timestamp 1666464484
transform 1 0 6999 0 1 10220
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_2
timestamp 1666464484
transform 1 0 6362 0 1 10011
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_3
timestamp 1666464484
transform 1 0 8417 0 1 10011
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_4
timestamp 1666464484
transform 1 0 7890 0 1 10428
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_5
timestamp 1666464484
transform 1 0 6072 0 1 10428
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_6
timestamp 1666464484
transform 1 0 4952 0 1 10637
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_7
timestamp 1666464484
transform 1 0 3937 0 1 10845
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_8
timestamp 1666464484
transform 1 0 1698 0 1 11262
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_9
timestamp 1666464484
transform 1 0 9524 0 1 10845
box 0 0 1 1
use M3_M2$$43371564_256x8m81  M3_M2$$43371564_256x8m81_10
timestamp 1666464484
transform 1 0 9537 0 1 11471
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_0
timestamp 1666464484
transform 1 0 6953 0 1 13665
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_1
timestamp 1666464484
transform 1 0 6505 0 1 13665
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_2
timestamp 1666464484
transform 1 0 8072 0 1 14006
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_3
timestamp 1666464484
transform 1 0 7625 0 1 14006
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_4
timestamp 1666464484
transform 1 0 9192 0 1 14346
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_5
timestamp 1666464484
transform 1 0 8744 0 1 14346
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_6
timestamp 1666464484
transform 1 0 905 0 1 11965
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_7
timestamp 1666464484
transform 1 0 1353 0 1 11965
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_8
timestamp 1666464484
transform 1 0 2473 0 1 12305
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_9
timestamp 1666464484
transform 1 0 2025 0 1 12305
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_10
timestamp 1666464484
transform 1 0 3593 0 1 12645
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_11
timestamp 1666464484
transform 1 0 3145 0 1 12645
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_12
timestamp 1666464484
transform 1 0 4713 0 1 12985
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_13
timestamp 1666464484
transform 1 0 4265 0 1 12985
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_14
timestamp 1666464484
transform 1 0 5833 0 1 13325
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_15
timestamp 1666464484
transform 1 0 5385 0 1 13325
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_16
timestamp 1666464484
transform -1 0 11432 0 -1 12305
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_17
timestamp 1666464484
transform -1 0 10984 0 -1 12305
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_18
timestamp 1666464484
transform -1 0 12552 0 -1 12645
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_19
timestamp 1666464484
transform -1 0 12104 0 -1 12645
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_20
timestamp 1666464484
transform -1 0 13672 0 -1 12985
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_21
timestamp 1666464484
transform -1 0 13224 0 -1 12985
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_22
timestamp 1666464484
transform -1 0 14792 0 -1 13325
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_23
timestamp 1666464484
transform -1 0 14344 0 -1 13325
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_24
timestamp 1666464484
transform -1 0 15912 0 -1 13665
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_25
timestamp 1666464484
transform -1 0 15464 0 -1 13665
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_26
timestamp 1666464484
transform -1 0 17032 0 -1 14006
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_27
timestamp 1666464484
transform -1 0 16584 0 -1 14006
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_28
timestamp 1666464484
transform -1 0 17704 0 -1 14346
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_29
timestamp 1666464484
transform -1 0 18152 0 -1 14346
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_30
timestamp 1666464484
transform 1 0 10086 0 1 11054
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_31
timestamp 1666464484
transform -1 0 10312 0 -1 11965
box 0 0 1 1
use M3_M2$$46895148_256x8m81  M3_M2$$46895148_256x8m81_32
timestamp 1666464484
transform -1 0 9864 0 -1 11965
box 0 0 1 1
use M3_M2$$47632428_256x8m81  M3_M2$$47632428_256x8m81_0
timestamp 1666464484
transform -1 0 10023 0 1 478
box -1962 -176 1962 176
use M3_M2$$47633452_256x8m81  M3_M2$$47633452_256x8m81_0
timestamp 1666464484
transform -1 0 10157 0 1 1313
box -1857 -176 1857 176
use nmos_1p2$$47342636_256x8m81  nmos_1p2$$47342636_256x8m81_0
timestamp 1666464484
transform -1 0 6441 0 1 997
box -119 -73 177 316
use nmos_5p04310590878160_256x8m81  nmos_5p04310590878160_256x8m81_0
timestamp 1666464484
transform -1 0 7842 0 1 1002
box -88 -44 208 426
use nmos_5p04310590878160_256x8m81  nmos_5p04310590878160_256x8m81_1
timestamp 1666464484
transform -1 0 8066 0 1 1002
box -88 -44 208 426
use pmos_1p2$$47109164_256x8m81  pmos_1p2$$47109164_256x8m81_0
timestamp 1666464484
transform -1 0 6559 0 1 281
box -239 -120 521 462
use ypredec1_bot_256x8m81  ypredec1_bot_256x8m81_0
timestamp 1666464484
transform 1 0 3766 0 1 1027
box -20 -633 1953 7883
use ypredec1_bot_256x8m81  ypredec1_bot_256x8m81_1
timestamp 1666464484
transform 1 0 384 0 1 1027
box -20 -633 1953 7883
use ypredec1_bot_256x8m81  ypredec1_bot_256x8m81_2
timestamp 1666464484
transform 1 0 2075 0 1 1027
box -20 -633 1953 7883
use ypredec1_xax8_256x8m81  ypredec1_xax8_256x8m81_0
timestamp 1666464484
transform 1 0 5624 0 1 1528
box -1 -55 6822 7396
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_0
timestamp 1666464484
transform 1 0 255 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_1
timestamp 1666464484
transform 1 0 1375 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_2
timestamp 1666464484
transform 1 0 2495 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_3
timestamp 1666464484
transform 1 0 3615 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_4
timestamp 1666464484
transform 1 0 4735 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_5
timestamp 1666464484
transform 1 0 5855 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_6
timestamp 1666464484
transform 1 0 6975 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_7
timestamp 1666464484
transform 1 0 10335 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_8
timestamp 1666464484
transform 1 0 11455 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_9
timestamp 1666464484
transform 1 0 12575 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_10
timestamp 1666464484
transform 1 0 13695 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_11
timestamp 1666464484
transform 1 0 14815 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_12
timestamp 1666464484
transform 1 0 15935 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_13
timestamp 1666464484
transform 1 0 17055 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_14
timestamp 1666464484
transform 1 0 9215 0 1 9054
box -1 -1 1931 7382
use ypredec1_ys_256x8m81  ypredec1_ys_256x8m81_15
timestamp 1666464484
transform 1 0 8095 0 1 9054
box -1 -1 1931 7382
<< labels >>
rlabel metal3 s 993 13665 993 13665 4 ly[5]
port 1 nsew
rlabel metal3 s 993 13325 993 13325 4 ly[4]
port 2 nsew
rlabel metal3 s 993 14346 993 14346 4 ly[7]
port 3 nsew
rlabel metal3 s 993 12985 993 12985 4 ly[3]
port 4 nsew
rlabel metal3 s 993 12645 993 12645 4 ly[2]
port 5 nsew
rlabel metal3 s 993 12305 993 12305 4 ly[1]
port 6 nsew
rlabel metal3 s 993 11965 993 11965 4 ly[0]
port 7 nsew
rlabel metal3 s 25537 11965 25537 11965 4 ry[0]
port 8 nsew
rlabel metal3 s 25537 12305 25537 12305 4 ry[1]
port 9 nsew
rlabel metal3 s 25537 12645 25537 12645 4 ry[2]
port 10 nsew
rlabel metal3 s 25537 12985 25537 12985 4 ry[3]
port 11 nsew
rlabel metal3 s 25537 13325 25537 13325 4 ry[4]
port 12 nsew
rlabel metal3 s 25537 13665 25537 13665 4 ry[5]
port 13 nsew
rlabel metal3 s 25537 14006 25537 14006 4 ry[6]
port 14 nsew
rlabel metal3 s 25537 14346 25537 14346 4 ry[7]
port 15 nsew
rlabel metal3 s 993 14006 993 14006 4 ly[6]
port 16 nsew
rlabel metal2 s 8314 855 8314 855 4 men
port 17 nsew
rlabel metal2 s 5257 673 5257 673 4 A[0]
port 18 nsew
rlabel metal2 s 3566 673 3566 673 4 A[1]
port 19 nsew
rlabel metal2 s 1875 673 1875 673 4 A[2]
port 20 nsew
rlabel metal2 s 7466 1335 7466 1335 4 clk
port 21 nsew
<< properties >>
string GDS_END 1827244
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1805738
<< end >>
