magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 1120 844
rect 242 582 310 724
rect 535 532 581 678
rect 728 582 796 724
rect 916 532 1032 678
rect 141 325 330 430
rect 535 442 1032 532
rect 141 122 203 325
rect 916 260 1032 442
rect 535 213 1032 260
rect 300 60 368 153
rect 535 114 581 213
rect 748 60 816 153
rect 916 114 1032 213
rect 0 -60 1120 60
<< obsm1 >>
rect 49 525 95 678
rect 49 478 426 525
rect 49 114 95 478
rect 380 378 426 478
rect 380 310 835 378
<< labels >>
rlabel metal1 s 141 325 330 430 6 I
port 1 nsew default input
rlabel metal1 s 141 122 203 325 6 I
port 1 nsew default input
rlabel metal1 s 916 532 1032 678 6 Z
port 2 nsew default output
rlabel metal1 s 535 532 581 678 6 Z
port 2 nsew default output
rlabel metal1 s 535 442 1032 532 6 Z
port 2 nsew default output
rlabel metal1 s 916 260 1032 442 6 Z
port 2 nsew default output
rlabel metal1 s 535 213 1032 260 6 Z
port 2 nsew default output
rlabel metal1 s 916 114 1032 213 6 Z
port 2 nsew default output
rlabel metal1 s 535 114 581 213 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 1120 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 728 582 796 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 242 582 310 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 748 60 816 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 300 60 368 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1120 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1312544
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1309260
<< end >>
