magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -1386 23 1386 77
rect -1386 -23 -1329 23
rect -1283 -23 -1166 23
rect -1120 -23 -1003 23
rect -957 -23 -839 23
rect -793 -23 -676 23
rect -630 -23 -513 23
rect -467 -23 -350 23
rect -304 -23 -186 23
rect -140 -23 -23 23
rect 23 -23 140 23
rect 186 -23 304 23
rect 350 -23 467 23
rect 513 -23 630 23
rect 676 -23 793 23
rect 839 -23 957 23
rect 1003 -23 1120 23
rect 1166 -23 1283 23
rect 1329 -23 1386 23
rect -1386 -78 1386 -23
<< psubdiffcont >>
rect -1329 -23 -1283 23
rect -1166 -23 -1120 23
rect -1003 -23 -957 23
rect -839 -23 -793 23
rect -676 -23 -630 23
rect -513 -23 -467 23
rect -350 -23 -304 23
rect -186 -23 -140 23
rect -23 -23 23 23
rect 140 -23 186 23
rect 304 -23 350 23
rect 467 -23 513 23
rect 630 -23 676 23
rect 793 -23 839 23
rect 957 -23 1003 23
rect 1120 -23 1166 23
rect 1283 -23 1329 23
<< metal1 >>
rect -254 57 1185 58
rect -1366 23 1366 57
rect -1366 -23 -1329 23
rect -1283 -23 -1166 23
rect -1120 -23 -1003 23
rect -957 -23 -839 23
rect -793 -23 -676 23
rect -630 -23 -513 23
rect -467 -23 -350 23
rect -304 -23 -186 23
rect -140 -23 -23 23
rect 23 -23 140 23
rect 186 -23 304 23
rect 350 -23 467 23
rect 513 -23 630 23
rect 676 -23 793 23
rect 839 -23 957 23
rect 1003 -23 1120 23
rect 1166 -23 1283 23
rect 1329 -23 1366 23
rect -1366 -58 1366 -23
<< properties >>
string GDS_END 949458
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 948126
<< end >>
