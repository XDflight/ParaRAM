magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -65 26 1751 67
rect -65 -26 -26 26
rect 26 -26 185 26
rect 237 -26 396 26
rect 448 -26 607 26
rect 659 -26 818 26
rect 870 -26 1028 26
rect 1080 -26 1239 26
rect 1291 -26 1450 26
rect 1502 -26 1661 26
rect 1713 -26 1751 26
rect -65 -192 1751 -26
rect -65 -244 -26 -192
rect 26 -244 185 -192
rect 237 -244 396 -192
rect 448 -244 607 -192
rect 659 -244 818 -192
rect 870 -244 1028 -192
rect 1080 -244 1239 -192
rect 1291 -244 1450 -192
rect 1502 -244 1661 -192
rect 1713 -244 1751 -192
rect -65 -409 1751 -244
rect -65 -461 -26 -409
rect 26 -461 185 -409
rect 237 -461 396 -409
rect 448 -461 607 -409
rect 659 -461 818 -409
rect 870 -461 1028 -409
rect 1080 -461 1239 -409
rect 1291 -461 1450 -409
rect 1502 -461 1661 -409
rect 1713 -461 1751 -409
rect -65 -502 1751 -461
<< via1 >>
rect -26 -26 26 26
rect 185 -26 237 26
rect 396 -26 448 26
rect 607 -26 659 26
rect 818 -26 870 26
rect 1028 -26 1080 26
rect 1239 -26 1291 26
rect 1450 -26 1502 26
rect 1661 -26 1713 26
rect -26 -244 26 -192
rect 185 -244 237 -192
rect 396 -244 448 -192
rect 607 -244 659 -192
rect 818 -244 870 -192
rect 1028 -244 1080 -192
rect 1239 -244 1291 -192
rect 1450 -244 1502 -192
rect 1661 -244 1713 -192
rect -26 -461 26 -409
rect 185 -461 237 -409
rect 396 -461 448 -409
rect 607 -461 659 -409
rect 818 -461 870 -409
rect 1028 -461 1080 -409
rect 1239 -461 1291 -409
rect 1450 -461 1502 -409
rect 1661 -461 1713 -409
<< metal2 >>
rect -64 26 1751 67
rect -64 -26 -26 26
rect 26 -26 185 26
rect 237 -26 396 26
rect 448 -26 607 26
rect 659 -26 818 26
rect 870 -26 1028 26
rect 1080 -26 1239 26
rect 1291 -26 1450 26
rect 1502 -26 1661 26
rect 1713 -26 1751 26
rect -64 -192 1751 -26
rect -64 -244 -26 -192
rect 26 -244 185 -192
rect 237 -244 396 -192
rect 448 -244 607 -192
rect 659 -244 818 -192
rect 870 -244 1028 -192
rect 1080 -244 1239 -192
rect 1291 -244 1450 -192
rect 1502 -244 1661 -192
rect 1713 -244 1751 -192
rect -64 -409 1751 -244
rect -64 -461 -26 -409
rect 26 -461 185 -409
rect 237 -461 396 -409
rect 448 -461 607 -409
rect 659 -461 818 -409
rect 870 -461 1028 -409
rect 1080 -461 1239 -409
rect 1291 -461 1450 -409
rect 1502 -461 1661 -409
rect 1713 -461 1751 -409
rect -64 -502 1751 -461
<< properties >>
string GDS_END 1663334
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1661474
<< end >>
