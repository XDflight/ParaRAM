magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -532 23867 21664 29129
rect -532 17407 21671 19961
<< mvpmos >>
rect 4103 27950 4223 28632
rect 4328 27950 4448 28632
rect 4794 27950 4914 28632
rect 5019 27950 5139 28632
rect 14903 27950 15023 28632
rect 15128 27950 15248 28632
rect 15594 27950 15714 28632
rect 15819 27950 15939 28632
rect 4103 27175 4223 27857
rect 4328 27175 4448 27857
rect 4794 27175 4914 27857
rect 5019 27175 5139 27857
rect 14903 27175 15023 27857
rect 15128 27175 15248 27857
rect 15594 27175 15714 27857
rect 15819 27175 15939 27857
<< mvpdiff >>
rect 3997 27950 4103 28632
rect 4223 27950 4328 28632
rect 4448 27950 4554 28632
rect 4688 27950 4794 28632
rect 4914 27950 5019 28632
rect 5139 27950 5245 28632
rect 14797 27950 14903 28632
rect 15023 27950 15128 28632
rect 15248 27950 15354 28632
rect 15488 27950 15594 28632
rect 15714 27950 15819 28632
rect 15939 27950 16045 28632
rect 3997 27175 4103 27857
rect 4223 27175 4328 27857
rect 4448 27175 4554 27857
rect 4688 27175 4794 27857
rect 4914 27175 5019 27857
rect 5139 27175 5245 27857
rect 14797 27175 14903 27857
rect 15023 27175 15128 27857
rect 15248 27175 15354 27857
rect 15488 27175 15594 27857
rect 15714 27175 15819 27857
rect 15939 27175 16045 27857
<< metal1 >>
rect -994 29890 -918 29900
rect -844 29890 -714 30180
rect -994 29888 640 29890
rect -994 29732 -982 29888
rect -930 29732 640 29888
rect 4539 29867 4703 30180
rect 9939 29900 10103 30180
rect 9791 29888 10103 29900
rect -994 29720 640 29732
rect 9791 29732 9803 29888
rect 9959 29867 10103 29888
rect 15339 29867 15503 30180
rect 20739 29900 20903 30180
rect 20739 29888 21000 29900
rect 20739 29867 20832 29888
rect 9959 29732 9971 29867
rect 9791 29720 9971 29732
rect 20820 29732 20832 29867
rect 20988 29732 21000 29888
rect 20820 29720 21000 29732
rect 14849 16092 15238 16230
rect 15664 16092 16243 16230
<< via1 >>
rect -982 29732 -930 29888
rect 9803 29732 9959 29888
rect 20832 29732 20988 29888
<< metal2 >>
rect -1009 29987 -909 31176
rect -1009 29931 -983 29987
rect -927 29931 -909 29987
rect -1009 29888 -909 29931
rect -1009 29855 -982 29888
rect -930 29855 -909 29888
rect -1009 29799 -983 29855
rect -927 29799 -909 29855
rect -1009 29732 -982 29799
rect -930 29732 -909 29799
rect -1009 29723 -909 29732
rect -1009 29667 -983 29723
rect -927 29667 -909 29723
rect -1009 29591 -909 29667
rect -1009 29535 -983 29591
rect -927 29535 -909 29591
rect -1009 27521 -909 29535
rect -827 29107 -738 29955
rect -827 29069 -733 29107
rect -827 29013 -808 29069
rect -752 29013 -733 29069
rect -827 28883 -733 29013
rect -827 28827 -808 28883
rect -752 28827 -733 28883
rect -827 28788 -733 28827
rect -827 21746 -738 28788
rect -649 27516 -549 31176
rect 9791 29987 9891 31176
rect 9791 29931 9814 29987
rect 9870 29931 9891 29987
rect 9791 29900 9891 29931
rect 9791 29888 9971 29900
rect 9791 29732 9803 29888
rect 9959 29732 9971 29888
rect 9791 29723 9971 29732
rect 9791 29667 9814 29723
rect 9870 29720 9971 29723
rect 9870 29667 9891 29720
rect 9791 29591 9891 29667
rect 9791 29535 9814 29591
rect 9870 29535 9891 29591
rect 9791 27540 9891 29535
rect 10151 27539 10251 31176
rect 20591 27524 20691 31176
rect 20951 29987 21051 31176
rect 20951 29931 20975 29987
rect 21031 29931 21051 29987
rect 20951 29900 21051 29931
rect 20820 29888 21051 29900
rect 20820 29732 20832 29888
rect 20988 29855 21051 29888
rect 21031 29799 21051 29855
rect 20988 29732 21051 29799
rect 20820 29723 21051 29732
rect 20820 29720 20975 29723
rect 20951 29667 20975 29720
rect 21031 29667 21051 29723
rect 20951 29591 21051 29667
rect 20951 29535 20975 29591
rect 21031 29535 21051 29591
rect 20951 27527 21051 29535
<< via2 >>
rect -983 29931 -927 29987
rect -983 29799 -982 29855
rect -982 29799 -930 29855
rect -930 29799 -927 29855
rect -983 29667 -927 29723
rect -983 29535 -927 29591
rect -808 29013 -752 29069
rect -808 28827 -752 28883
rect 9814 29931 9870 29987
rect 9814 29799 9870 29855
rect 9814 29667 9870 29723
rect 9814 29535 9870 29591
rect 20975 29931 21031 29987
rect 20975 29799 20988 29855
rect 20988 29799 21031 29855
rect 20975 29667 21031 29723
rect 20975 29535 21031 29591
<< metal3 >>
rect -1115 38517 22810 38877
rect -1115 37737 22810 38097
rect -1115 36717 22810 37077
rect -1115 35937 22810 36297
rect -1115 34917 22810 35277
rect -1115 34137 22810 34497
rect -1115 33117 22810 33477
rect -1115 32337 22810 32697
rect -1115 31317 22810 31677
rect -1115 30537 22810 30897
rect -1186 29987 22164 29997
rect -1186 29931 -983 29987
rect -927 29931 9814 29987
rect 9870 29931 20975 29987
rect 21031 29931 22164 29987
rect -1186 29855 22164 29931
rect -1186 29799 -983 29855
rect -927 29799 9814 29855
rect 9870 29799 20975 29855
rect 21031 29799 22164 29855
rect -1186 29723 22164 29799
rect -1186 29667 -983 29723
rect -927 29667 9814 29723
rect 9870 29667 20975 29723
rect 21031 29667 22164 29723
rect -1186 29591 22164 29667
rect -1186 29535 -983 29591
rect -927 29535 9814 29591
rect 9870 29535 20975 29591
rect 21031 29535 22164 29591
rect -1186 29517 22164 29535
rect -826 29106 -733 29107
rect -1186 29069 22164 29106
rect -1186 29013 -808 29069
rect -752 29013 22164 29069
rect -1186 28883 22164 29013
rect -1186 28827 -808 28883
rect -752 28827 22164 28883
rect -1186 27297 22164 28827
rect -672 21090 21329 21305
rect -672 20768 21329 20983
rect -672 20447 21329 20662
rect -672 20125 21329 20340
rect -672 19433 21329 19648
rect -672 19111 21329 19326
rect -672 18790 21329 19005
rect -672 18468 21329 18683
rect -672 17919 21329 18361
rect -672 16808 21329 17263
rect -672 12997 21329 15720
rect -672 11578 20757 12711
rect -672 9309 21329 11578
rect -701 8442 21329 9159
rect 20900 7827 21329 7828
rect -701 7017 21329 7827
rect -672 5155 21329 6472
rect -672 4929 20872 5005
rect -672 3134 21329 4496
rect -672 1961 21329 2576
rect -672 1285 21329 1854
rect -672 747 21329 1179
rect -672 155 21329 610
rect -709 -959 21420 -504
rect -709 -1598 21420 -1247
rect -709 -1810 21420 -1722
rect -709 -2041 21420 -1953
rect -709 -2517 21420 -2166
rect -709 -3242 21420 -2787
use M2_M1431058998329_64x8m81  M2_M1431058998329_64x8m81_0
timestamp 1666464484
transform 1 0 -956 0 1 29810
box 0 0 1 1
use M2_M143105899832112_64x8m81  M2_M143105899832112_64x8m81_0
timestamp 1666464484
transform 1 0 9881 0 1 29810
box 0 0 1 1
use M2_M143105899832112_64x8m81  M2_M143105899832112_64x8m81_1
timestamp 1666464484
transform 1 0 20910 0 1 29810
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_0
timestamp 1666464484
transform 1 0 9842 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_1
timestamp 1666464484
transform 1 0 -955 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_2
timestamp 1666464484
transform 1 0 21003 0 1 29761
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_0
timestamp 1666464484
transform 1 0 20640 0 1 28318
box -38 -764 38 764
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_1
timestamp 1666464484
transform 1 0 -598 0 1 28318
box -38 -764 38 764
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_2
timestamp 1666464484
transform 1 0 10205 0 1 28318
box -38 -764 38 764
use col_64a_64x8m81_0  col_64a_64x8m81_0_0
timestamp 1666464484
transform 1 0 -1079 0 1 31107
box -68 -68 22268 7268
use dcap_103_novia_64x8m81  dcap_103_novia_64x8m81_0
array 0 35 619 0 0 0
timestamp 1666464484
transform 1 0 -827 0 1 29009
box -203 -284 822 881
use ldummy_64x4_64x8m81  ldummy_64x4_64x8m81_0
timestamp 1666464484
transform 1 0 -541 0 1 30030
box -636 76 22573 9277
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_0
timestamp 1666464484
transform -1 0 21008 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_1
timestamp 1666464484
transform -1 0 10208 0 1 6
box -269 -3400 7633 31133
use saout_m2_64x8m81  saout_m2_64x8m81_0
timestamp 1666464484
transform 1 0 -966 0 1 -1
box -269 -3393 7633 31140
use saout_m2_64x8m81  saout_m2_64x8m81_1
timestamp 1666464484
transform 1 0 9834 0 1 -1
box -269 -3393 7633 31140
use via2_x2_64x8m81  via2_x2_64x8m81_0
timestamp 1666464484
transform 1 0 -826 0 1 28789
box 0 0 1 1
<< labels >>
rlabel metal1 s 5690 15928 5690 15928 4 pcb[2]
port 1 nsew
rlabel metal1 s 3660 15928 3660 15928 4 pcb[3]
port 2 nsew
rlabel metal1 s 16496 15928 16496 15928 4 pcb[0]
port 3 nsew
rlabel metal1 s 14155 15928 14155 15928 4 pcb[1]
port 4 nsew
rlabel metal1 s 920 18163 920 18163 4 vdd
port 5 nsew
flabel metal1 s -808 31106 -808 31106 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal1 s -367 -3355 -367 -3355 0 FreeSans 600 0 0 0 WEN[3]
port 7 nsew
flabel metal1 s 9597 -3329 9597 -3329 0 FreeSans 600 0 0 0 WEN[2]
port 8 nsew
flabel metal1 s 10395 -3329 10395 -3329 0 FreeSans 600 0 0 0 WEN[1]
port 9 nsew
flabel metal1 s 20398 -3329 20398 -3329 0 FreeSans 600 0 0 0 WEN[0]
port 10 nsew
rlabel metal1 s 16437 15928 16437 15928 4 pcb[0]
port 3 nsew
rlabel metal1 s 14224 15928 14224 15928 4 pcb[1]
port 4 nsew
rlabel metal1 s 3672 15928 3672 15928 4 pcb[3]
port 2 nsew
rlabel metal1 s 5615 15928 5615 15928 4 pcb[2]
port 1 nsew
flabel metal1 s -367 -3355 -367 -3355 0 FreeSans 600 0 0 0 WEN[3]
port 7 nsew
flabel metal1 s 9740 -3329 9740 -3329 0 FreeSans 600 0 0 0 WEN[2]
port 8 nsew
flabel metal1 s 10394 -3329 10394 -3329 0 FreeSans 600 0 0 0 WEN[1]
port 9 nsew
flabel metal1 s 20462 -3329 20462 -3329 0 FreeSans 600 0 0 0 WEN[0]
port 10 nsew
rlabel metal3 s 701 37868 701 37868 4 WL[7]
port 11 nsew
rlabel metal3 s 701 36968 701 36968 4 WL[6]
port 12 nsew
rlabel metal3 s 701 36068 701 36068 4 WL[5]
port 13 nsew
rlabel metal3 s 701 35168 701 35168 4 WL[4]
port 14 nsew
rlabel metal3 s 701 34268 701 34268 4 WL[3]
port 15 nsew
rlabel metal3 s 701 33368 701 33368 4 WL[2]
port 16 nsew
rlabel metal3 s 701 32468 701 32468 4 WL[1]
port 17 nsew
rlabel metal3 s 701 31568 701 31568 4 WL[0]
port 18 nsew
rlabel metal3 s 870 1467 870 1467 4 men
port 19 nsew
rlabel metal3 s 797 18592 797 18592 4 ypass[0]
port 20 nsew
rlabel metal3 s 797 18914 797 18914 4 ypass[1]
port 21 nsew
rlabel metal3 s 797 19231 797 19231 4 ypass[2]
port 22 nsew
rlabel metal3 s 797 19548 797 19548 4 ypass[3]
port 23 nsew
rlabel metal3 s 797 20204 797 20204 4 ypass[4]
port 24 nsew
rlabel metal3 s 797 20528 797 20528 4 ypass[5]
port 25 nsew
rlabel metal3 s 797 20845 797 20845 4 ypass[6]
port 26 nsew
rlabel metal3 s 797 21162 797 21162 4 ypass[7]
port 27 nsew
rlabel metal3 s 867 1467 867 1467 4 men
port 19 nsew
flabel metal3 s -334 8814 -334 8814 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 386 -334 386 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -305 1002 -305 1002 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 2322 -305 2322 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 5923 -305 5923 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 11468 -305 11468 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 22970 -305 22970 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 29782 -305 29782 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -334 3858 -334 3858 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 7580 -334 7580 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 14009 -334 14009 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 18141 -334 18141 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 27925 -334 27925 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 -708 -334 -708 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -334 -3027 -334 -3027 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -305 -1478 -305 -1478 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -305 -2341 -305 -2341 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s 793 -1999 793 -1999 0 FreeSans 2000 0 0 0 GWEN
port 29 nsew
flabel metal3 s -325 4973 -325 4973 0 FreeSans 2000 0 0 0 GWE
port 30 nsew
rlabel metal3 s -728 34270 -728 34270 4 WL[3]
port 15 nsew
rlabel metal3 s 797 18591 797 18591 4 ypass[0]
port 20 nsew
rlabel metal3 s 797 18913 797 18913 4 ypass[1]
port 21 nsew
rlabel metal3 s 797 19548 797 19548 4 ypass[3]
port 23 nsew
rlabel metal3 s 797 20203 797 20203 4 ypass[4]
port 24 nsew
rlabel metal3 s 797 20527 797 20527 4 ypass[5]
port 25 nsew
rlabel metal3 s 797 21162 797 21162 4 ypass[7]
port 27 nsew
rlabel metal3 s 868 1466 868 1466 4 men
port 19 nsew
flabel metal3 s -327 4977 -327 4977 0 FreeSans 2000 0 0 0 GWE
port 30 nsew
flabel metal3 s -327 -3052 -327 -3052 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 -738 -327 -738 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
rlabel metal3 s -728 33370 -728 33370 4 WL[2]
port 16 nsew
rlabel metal3 s -728 32470 -728 32470 4 WL[1]
port 17 nsew
flabel metal3 s -327 390 -327 390 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
rlabel metal3 s -728 37870 -728 37870 4 WL[7]
port 11 nsew
rlabel metal3 s -728 36970 -728 36970 4 WL[6]
port 12 nsew
rlabel metal3 s -728 36070 -728 36070 4 WL[5]
port 13 nsew
rlabel metal3 s -728 35170 -728 35170 4 WL[4]
port 14 nsew
rlabel metal3 s -728 31570 -728 31570 4 WL[0]
port 18 nsew
rlabel metal3 s 798 20844 798 20844 4 ypass[6]
port 26 nsew
rlabel metal3 s 798 19230 798 19230 4 ypass[2]
port 22 nsew
flabel metal3 s -327 998 -327 998 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 2325 -327 2325 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 3859 -327 3859 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 7582 -327 7582 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 14010 -327 14010 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 18137 -327 18137 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 27926 -327 27926 0 FreeSans 2000 0 0 0 VDD
port 6 nsew
flabel metal3 s -327 29771 -327 29771 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 22970 -327 22970 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 11464 -327 11464 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
flabel metal3 s -327 5924 -327 5924 0 FreeSans 2000 0 0 0 VSS
port 28 nsew
rlabel metal2 s -454 104 -454 104 4 din[0]
port 31 nsew
rlabel metal2 s 9695 104 9695 104 4 din[1]
port 32 nsew
rlabel metal2 s 10331 104 10331 104 4 din[2]
port 33 nsew
rlabel metal2 s 8835 104 8835 104 4 q[1]
port 34 nsew
rlabel metal2 s 19234 29015 19234 29015 4 b[1]
port 35 nsew
rlabel metal2 s 17793 29015 17793 29015 4 b[4]
port 36 nsew
rlabel metal2 s 15518 29015 15518 29015 4 b[7]
port 37 nsew
rlabel metal2 s 14077 29015 14077 29015 4 b[10]
port 38 nsew
rlabel metal2 s 11802 29015 11802 29015 4 b[13]
port 39 nsew
rlabel metal2 s 9466 29015 9466 29015 4 b[16]
port 40 nsew
rlabel metal2 s 7190 29015 7190 29015 4 b[19]
port 41 nsew
rlabel metal2 s 5750 29015 5750 29015 4 b[22]
port 42 nsew
rlabel metal2 s 3475 29015 3475 29015 4 b[25]
port 43 nsew
rlabel metal2 s 2034 29015 2034 29015 4 b[28]
port 44 nsew
rlabel metal2 s -241 29015 -241 29015 4 b[31]
port 45 nsew
rlabel metal2 s 20495 104 20495 104 4 din[3]
port 46 nsew
rlabel metal2 s 382 104 382 104 4 q[0]
port 47 nsew
rlabel metal2 s 11187 104 11187 104 4 q[2]
port 48 nsew
rlabel metal2 s 19655 104 19655 104 4 q[3]
port 49 nsew
rlabel metal2 s 998 29015 998 29015 4 b[29]
port 50 nsew
rlabel metal2 s 3273 29015 3273 29015 4 b[26]
port 51 nsew
rlabel metal2 s 4713 29015 4713 29015 4 b[23]
port 52 nsew
rlabel metal2 s 6988 29015 6988 29015 4 b[20]
port 53 nsew
rlabel metal2 s 8429 29015 8429 29015 4 b[17]
port 54 nsew
rlabel metal2 s 11600 29015 11600 29015 4 b[14]
port 55 nsew
rlabel metal2 s 13041 29015 13041 29015 4 b[11]
port 56 nsew
rlabel metal2 s 15316 29015 15316 29015 4 b[8]
port 57 nsew
rlabel metal2 s 16757 29015 16757 29015 4 b[5]
port 58 nsew
rlabel metal2 s 19032 29015 19032 29015 4 b[2]
port 59 nsew
rlabel metal2 s 19853 29015 19853 29015 4 bb[0]
port 60 nsew
rlabel metal2 s 19651 29015 19651 29015 4 bb[1]
port 61 nsew
rlabel metal2 s 18614 29015 18614 29015 4 bb[2]
port 62 nsew
rlabel metal2 s 18412 29015 18412 29015 4 bb[3]
port 63 nsew
rlabel metal2 s 17376 29015 17376 29015 4 bb[4]
port 64 nsew
rlabel metal2 s 17174 29015 17174 29015 4 bb[5]
port 65 nsew
rlabel metal2 s 16137 29015 16137 29015 4 bb[6]
port 66 nsew
rlabel metal2 s 15935 29015 15935 29015 4 bb[7]
port 67 nsew
rlabel metal2 s 14899 29015 14899 29015 4 bb[8]
port 68 nsew
rlabel metal2 s 14697 29015 14697 29015 4 bb[9]
port 69 nsew
rlabel metal2 s 13660 29015 13660 29015 4 bb[10]
port 70 nsew
rlabel metal2 s 13458 29015 13458 29015 4 bb[11]
port 71 nsew
rlabel metal2 s 12422 29015 12422 29015 4 bb[12]
port 72 nsew
rlabel metal2 s 12220 29015 12220 29015 4 bb[13]
port 73 nsew
rlabel metal2 s 11183 29015 11183 29015 4 bb[14]
port 74 nsew
rlabel metal2 s 10981 29015 10981 29015 4 bb[15]
port 75 nsew
rlabel metal2 s 9048 29015 9048 29015 4 bb[16]
port 76 nsew
rlabel metal2 s 8846 29015 8846 29015 4 bb[17]
port 77 nsew
rlabel metal2 s 7810 29015 7810 29015 4 bb[18]
port 78 nsew
rlabel metal2 s 7608 29015 7608 29015 4 bb[19]
port 79 nsew
rlabel metal2 s 6571 29015 6571 29015 4 bb[20]
port 80 nsew
rlabel metal2 s 6369 29015 6369 29015 4 bb[21]
port 81 nsew
rlabel metal2 s 5333 29015 5333 29015 4 bb[22]
port 82 nsew
rlabel metal2 s 5131 29015 5131 29015 4 bb[23]
port 83 nsew
rlabel metal2 s 4094 29015 4094 29015 4 bb[24]
port 84 nsew
rlabel metal2 s 3892 29015 3892 29015 4 bb[25]
port 85 nsew
rlabel metal2 s 2856 29015 2856 29015 4 bb[26]
port 86 nsew
rlabel metal2 s 2654 29015 2654 29015 4 bb[27]
port 87 nsew
rlabel metal2 s 1617 29015 1617 29015 4 bb[28]
port 88 nsew
rlabel metal2 s 1415 29015 1415 29015 4 bb[29]
port 89 nsew
rlabel metal2 s 378 29015 378 29015 4 bb[30]
port 90 nsew
rlabel metal2 s 176 29015 176 29015 4 bb[31]
port 91 nsew
rlabel metal2 s 796 29015 796 29015 4 b[30]
port 92 nsew
rlabel metal2 s 2236 29015 2236 29015 4 b[27]
port 93 nsew
rlabel metal2 s 4511 29015 4511 29015 4 b[24]
port 94 nsew
rlabel metal2 s 10564 29015 10564 29015 4 b[15]
port 95 nsew
rlabel metal2 s 12839 29015 12839 29015 4 b[12]
port 96 nsew
rlabel metal2 s 14279 29015 14279 29015 4 b[9]
port 97 nsew
rlabel metal2 s 5952 29015 5952 29015 4 b[21]
port 98 nsew
rlabel metal2 s 20270 29015 20270 29015 4 b[0]
port 99 nsew
rlabel metal2 s 17995 29015 17995 29015 4 b[3]
port 100 nsew
rlabel metal2 s 16555 29015 16555 29015 4 b[6]
port 101 nsew
rlabel metal2 s 8227 29015 8227 29015 4 b[18]
port 102 nsew
rlabel metal3 701 38768 701 38768 4 WL[8]
rlabel metal3 -728 38770 -728 38770 4 WL[8]
<< properties >>
string FIXED_BBOX 15366 28635 15476 31202
string GDS_END 1646910
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1632686
string path 50.110 134.975 50.110 189.995 
<< end >>
