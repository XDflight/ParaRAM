magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 1448 574
<< mvpmos >>
rect 0 0 120 454
rect 224 0 344 454
rect 448 0 568 454
rect 672 0 792 454
rect 896 0 1016 454
rect 1120 0 1240 454
<< mvpdiff >>
rect -88 441 0 454
rect -88 395 -75 441
rect -29 395 0 441
rect -88 314 0 395
rect -88 268 -75 314
rect -29 268 0 314
rect -88 187 0 268
rect -88 141 -75 187
rect -29 141 0 187
rect -88 59 0 141
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 441 224 454
rect 120 395 149 441
rect 195 395 224 441
rect 120 314 224 395
rect 120 268 149 314
rect 195 268 224 314
rect 120 187 224 268
rect 120 141 149 187
rect 195 141 224 187
rect 120 59 224 141
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 441 448 454
rect 344 395 373 441
rect 419 395 448 441
rect 344 314 448 395
rect 344 268 373 314
rect 419 268 448 314
rect 344 187 448 268
rect 344 141 373 187
rect 419 141 448 187
rect 344 59 448 141
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 441 672 454
rect 568 395 597 441
rect 643 395 672 441
rect 568 314 672 395
rect 568 268 597 314
rect 643 268 672 314
rect 568 187 672 268
rect 568 141 597 187
rect 643 141 672 187
rect 568 59 672 141
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 441 896 454
rect 792 395 821 441
rect 867 395 896 441
rect 792 314 896 395
rect 792 268 821 314
rect 867 268 896 314
rect 792 187 896 268
rect 792 141 821 187
rect 867 141 896 187
rect 792 59 896 141
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 441 1120 454
rect 1016 395 1045 441
rect 1091 395 1120 441
rect 1016 314 1120 395
rect 1016 268 1045 314
rect 1091 268 1120 314
rect 1016 187 1120 268
rect 1016 141 1045 187
rect 1091 141 1120 187
rect 1016 59 1120 141
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 441 1328 454
rect 1240 395 1269 441
rect 1315 395 1328 441
rect 1240 314 1328 395
rect 1240 268 1269 314
rect 1315 268 1328 314
rect 1240 187 1328 268
rect 1240 141 1269 187
rect 1315 141 1328 187
rect 1240 59 1328 141
rect 1240 13 1269 59
rect 1315 13 1328 59
rect 1240 0 1328 13
<< mvpdiffc >>
rect -75 395 -29 441
rect -75 268 -29 314
rect -75 141 -29 187
rect -75 13 -29 59
rect 149 395 195 441
rect 149 268 195 314
rect 149 141 195 187
rect 149 13 195 59
rect 373 395 419 441
rect 373 268 419 314
rect 373 141 419 187
rect 373 13 419 59
rect 597 395 643 441
rect 597 268 643 314
rect 597 141 643 187
rect 597 13 643 59
rect 821 395 867 441
rect 821 268 867 314
rect 821 141 867 187
rect 821 13 867 59
rect 1045 395 1091 441
rect 1045 268 1091 314
rect 1045 141 1091 187
rect 1045 13 1091 59
rect 1269 395 1315 441
rect 1269 268 1315 314
rect 1269 141 1315 187
rect 1269 13 1315 59
<< polysilicon >>
rect 0 454 120 498
rect 224 454 344 498
rect 448 454 568 498
rect 672 454 792 498
rect 896 454 1016 498
rect 1120 454 1240 498
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
<< metal1 >>
rect -75 441 -29 454
rect -75 314 -29 395
rect -75 187 -29 268
rect -75 59 -29 141
rect -75 0 -29 13
rect 149 441 195 454
rect 149 314 195 395
rect 149 187 195 268
rect 149 59 195 141
rect 149 0 195 13
rect 373 441 419 454
rect 373 314 419 395
rect 373 187 419 268
rect 373 59 419 141
rect 373 0 419 13
rect 597 441 643 454
rect 597 314 643 395
rect 597 187 643 268
rect 597 59 643 141
rect 597 0 643 13
rect 821 441 867 454
rect 821 314 867 395
rect 821 187 867 268
rect 821 59 867 141
rect 821 0 867 13
rect 1045 441 1091 454
rect 1045 314 1091 395
rect 1045 187 1091 268
rect 1045 59 1091 141
rect 1045 0 1091 13
rect 1269 441 1315 454
rect 1269 314 1315 395
rect 1269 187 1315 268
rect 1269 59 1315 141
rect 1269 0 1315 13
<< labels >>
flabel metal1 s -52 227 -52 227 0 FreeSans 400 0 0 0 S
flabel metal1 s 1292 227 1292 227 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 227 172 227 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 227 396 227 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 227 620 227 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 227 844 227 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 227 1068 227 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 76824
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 72162
<< end >>
