magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 3894 870
<< pwell >>
rect -86 -86 3894 352
<< mvnmos >>
rect 124 156 244 232
rect 348 156 468 232
rect 660 156 780 232
rect 884 156 1004 232
rect 1108 156 1228 232
rect 1332 156 1452 232
rect 1784 156 1904 229
rect 2027 156 2147 229
rect 2424 156 2544 229
rect 2648 156 2768 229
rect 2872 156 2992 229
rect 3096 156 3216 229
rect 3320 156 3440 229
rect 3544 156 3664 229
<< mvpmos >>
rect 124 472 224 628
rect 424 472 524 628
rect 628 472 728 628
rect 884 472 984 628
rect 1108 472 1208 628
rect 1352 472 1452 628
rect 1772 509 1872 628
rect 2048 509 2148 628
rect 2444 509 2544 628
rect 2668 509 2768 628
rect 2872 509 2972 628
rect 3076 509 3176 628
rect 3320 509 3420 628
rect 3544 509 3644 628
<< mvndiff >>
rect 36 215 124 232
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 232
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 215 660 232
rect 468 169 525 215
rect 571 169 660 215
rect 468 156 660 169
rect 780 215 884 232
rect 780 169 809 215
rect 855 169 884 215
rect 780 156 884 169
rect 1004 215 1108 232
rect 1004 169 1033 215
rect 1079 169 1108 215
rect 1004 156 1108 169
rect 1228 215 1332 232
rect 1228 169 1257 215
rect 1303 169 1332 215
rect 1228 156 1332 169
rect 1452 215 1540 232
rect 1452 169 1481 215
rect 1527 169 1540 215
rect 1452 156 1540 169
rect 1634 215 1784 229
rect 1634 169 1647 215
rect 1693 169 1784 215
rect 1634 156 1784 169
rect 1904 215 2027 229
rect 1904 169 1933 215
rect 1979 169 2027 215
rect 1904 156 2027 169
rect 2147 215 2236 229
rect 2147 169 2177 215
rect 2223 169 2236 215
rect 2147 156 2236 169
rect 2336 216 2424 229
rect 2336 170 2349 216
rect 2395 170 2424 216
rect 2336 156 2424 170
rect 2544 216 2648 229
rect 2544 170 2573 216
rect 2619 170 2648 216
rect 2544 156 2648 170
rect 2768 216 2872 229
rect 2768 170 2797 216
rect 2843 170 2872 216
rect 2768 156 2872 170
rect 2992 216 3096 229
rect 2992 170 3021 216
rect 3067 170 3096 216
rect 2992 156 3096 170
rect 3216 216 3320 229
rect 3216 170 3245 216
rect 3291 170 3320 216
rect 3216 156 3320 170
rect 3440 216 3544 229
rect 3440 170 3469 216
rect 3515 170 3544 216
rect 3440 156 3544 170
rect 3664 216 3752 229
rect 3664 170 3693 216
rect 3739 170 3752 216
rect 3664 156 3752 170
<< mvpdiff >>
rect 36 579 124 628
rect 36 533 49 579
rect 95 533 124 579
rect 36 472 124 533
rect 224 579 424 628
rect 224 533 253 579
rect 299 533 424 579
rect 224 472 424 533
rect 524 605 628 628
rect 524 559 553 605
rect 599 559 628 605
rect 524 472 628 559
rect 728 574 884 628
rect 728 528 797 574
rect 843 528 884 574
rect 728 472 884 528
rect 984 615 1108 628
rect 984 569 1013 615
rect 1059 569 1108 615
rect 984 472 1108 569
rect 1208 571 1352 628
rect 1208 525 1257 571
rect 1303 525 1352 571
rect 1208 472 1352 525
rect 1452 571 1540 628
rect 1452 525 1481 571
rect 1527 525 1540 571
rect 1452 472 1540 525
rect 1637 590 1772 628
rect 1637 544 1650 590
rect 1696 544 1772 590
rect 1637 509 1772 544
rect 1872 590 2048 628
rect 1872 544 1919 590
rect 1965 544 2048 590
rect 1872 509 2048 544
rect 2148 590 2236 628
rect 2148 544 2177 590
rect 2223 544 2236 590
rect 2148 509 2236 544
rect 2356 574 2444 628
rect 2356 528 2369 574
rect 2415 528 2444 574
rect 2356 509 2444 528
rect 2544 615 2668 628
rect 2544 569 2593 615
rect 2639 569 2668 615
rect 2544 509 2668 569
rect 2768 574 2872 628
rect 2768 528 2797 574
rect 2843 528 2872 574
rect 2768 509 2872 528
rect 2972 574 3076 628
rect 2972 528 3001 574
rect 3047 528 3076 574
rect 2972 509 3076 528
rect 3176 609 3320 628
rect 3176 563 3228 609
rect 3274 563 3320 609
rect 3176 509 3320 563
rect 3420 609 3544 628
rect 3420 563 3449 609
rect 3495 563 3544 609
rect 3420 509 3544 563
rect 3644 609 3732 628
rect 3644 563 3673 609
rect 3719 563 3732 609
rect 3644 509 3732 563
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 525 169 571 215
rect 809 169 855 215
rect 1033 169 1079 215
rect 1257 169 1303 215
rect 1481 169 1527 215
rect 1647 169 1693 215
rect 1933 169 1979 215
rect 2177 169 2223 215
rect 2349 170 2395 216
rect 2573 170 2619 216
rect 2797 170 2843 216
rect 3021 170 3067 216
rect 3245 170 3291 216
rect 3469 170 3515 216
rect 3693 170 3739 216
<< mvpdiffc >>
rect 49 533 95 579
rect 253 533 299 579
rect 553 559 599 605
rect 797 528 843 574
rect 1013 569 1059 615
rect 1257 525 1303 571
rect 1481 525 1527 571
rect 1650 544 1696 590
rect 1919 544 1965 590
rect 2177 544 2223 590
rect 2369 528 2415 574
rect 2593 569 2639 615
rect 2797 528 2843 574
rect 3001 528 3047 574
rect 3228 563 3274 609
rect 3449 563 3495 609
rect 3673 563 3719 609
<< polysilicon >>
rect 628 720 2972 760
rect 124 628 224 672
rect 424 628 524 672
rect 628 628 728 720
rect 884 628 984 672
rect 1108 628 1208 672
rect 1352 628 1452 672
rect 1772 628 1872 672
rect 2048 628 2148 672
rect 2444 628 2544 672
rect 2668 628 2768 672
rect 2872 628 2972 720
rect 3076 720 3644 760
rect 3076 628 3176 720
rect 3320 628 3420 672
rect 3544 628 3644 720
rect 124 394 224 472
rect 124 348 141 394
rect 187 380 224 394
rect 424 439 524 472
rect 424 393 451 439
rect 497 393 524 439
rect 628 412 728 472
rect 424 380 524 393
rect 187 348 244 380
rect 124 232 244 348
rect 572 372 728 412
rect 884 408 984 472
rect 884 394 1004 408
rect 572 332 612 372
rect 348 292 612 332
rect 884 348 928 394
rect 974 348 1004 394
rect 660 311 780 324
rect 348 232 468 292
rect 660 265 679 311
rect 725 265 780 311
rect 660 232 780 265
rect 884 232 1004 348
rect 1108 364 1208 472
rect 1352 364 1452 472
rect 1772 409 1872 509
rect 2048 468 2148 509
rect 2048 422 2061 468
rect 2107 449 2148 468
rect 2444 449 2544 509
rect 2107 422 2544 449
rect 2668 426 2768 509
rect 2048 409 2544 422
rect 1772 369 2000 409
rect 1108 351 1724 364
rect 1108 305 1665 351
rect 1711 305 1724 351
rect 1952 361 2000 369
rect 1952 348 2329 361
rect 1952 321 2270 348
rect 1108 304 1724 305
rect 1108 232 1228 304
rect 1332 292 1724 304
rect 1784 308 1904 321
rect 1332 232 1452 292
rect 1784 262 1845 308
rect 1891 262 1904 308
rect 1784 229 1904 262
rect 2027 302 2270 321
rect 2316 302 2329 348
rect 2027 289 2329 302
rect 2027 229 2147 289
rect 2424 229 2544 409
rect 2648 414 2768 426
rect 2648 368 2682 414
rect 2728 368 2768 414
rect 2648 229 2768 368
rect 2872 405 2972 509
rect 3076 465 3176 509
rect 3320 431 3420 509
rect 3320 412 3440 431
rect 2872 392 3264 405
rect 2872 352 3205 392
rect 3096 346 3205 352
rect 3251 346 3264 392
rect 3096 333 3264 346
rect 3320 366 3353 412
rect 3399 366 3440 412
rect 2872 229 2992 273
rect 3096 229 3216 333
rect 3320 229 3440 366
rect 3544 355 3644 509
rect 3544 229 3664 355
rect 124 112 244 156
rect 348 112 468 156
rect 660 64 780 156
rect 884 112 1004 156
rect 1108 112 1228 156
rect 1332 112 1452 156
rect 1784 112 1904 156
rect 2027 112 2147 156
rect 2424 112 2544 156
rect 2648 112 2768 156
rect 2872 64 2992 156
rect 3096 112 3216 156
rect 3320 112 3440 156
rect 3544 64 3664 156
rect 660 24 3664 64
<< polycontact >>
rect 141 348 187 394
rect 451 393 497 439
rect 928 348 974 394
rect 679 265 725 311
rect 2061 422 2107 468
rect 1665 305 1711 351
rect 1845 262 1891 308
rect 2270 302 2316 348
rect 2682 368 2728 414
rect 3205 346 3251 392
rect 3353 366 3399 412
<< metal1 >>
rect 0 724 3808 844
rect 49 579 95 724
rect 542 620 947 666
rect 542 605 610 620
rect 542 594 553 605
rect 49 515 95 533
rect 141 394 202 590
rect 187 348 202 394
rect 49 215 95 226
rect 141 194 202 348
rect 252 579 299 590
rect 252 533 253 579
rect 252 215 299 533
rect 345 559 553 594
rect 599 559 610 605
rect 345 548 610 559
rect 345 314 391 548
rect 786 528 797 574
rect 843 528 855 574
rect 451 439 740 450
rect 497 393 740 439
rect 451 360 740 393
rect 345 268 458 314
rect 408 215 458 268
rect 660 311 740 360
rect 660 265 679 311
rect 725 265 740 311
rect 660 248 740 265
rect 786 215 855 528
rect 901 523 947 620
rect 1002 615 1070 724
rect 1002 569 1013 615
rect 1059 569 1070 615
rect 1134 631 1419 678
rect 1134 523 1180 631
rect 901 476 1180 523
rect 1246 525 1257 571
rect 1303 525 1320 571
rect 252 169 273 215
rect 319 169 330 215
rect 408 169 525 215
rect 571 169 582 215
rect 786 169 809 215
rect 49 60 95 169
rect 786 156 855 169
rect 901 394 1151 430
rect 901 348 928 394
rect 974 360 1151 394
rect 974 348 987 360
rect 901 110 987 348
rect 1033 215 1079 232
rect 1033 60 1079 169
rect 1246 215 1320 525
rect 1373 455 1419 631
rect 1481 571 1527 724
rect 1481 514 1527 525
rect 1573 590 1696 601
rect 1573 544 1650 590
rect 1573 533 1696 544
rect 1742 544 1919 590
rect 1965 544 1976 590
rect 1573 455 1619 533
rect 1373 409 1619 455
rect 1246 169 1257 215
rect 1303 169 1320 215
rect 1246 120 1320 169
rect 1481 215 1527 232
rect 1481 60 1527 169
rect 1573 226 1619 409
rect 1742 364 1788 544
rect 2033 468 2107 664
rect 2033 430 2061 468
rect 1665 351 1788 364
rect 1711 305 1788 351
rect 1665 292 1788 305
rect 1573 215 1696 226
rect 1573 169 1647 215
rect 1693 169 1696 215
rect 1742 215 1788 292
rect 1834 422 2061 430
rect 1834 354 2107 422
rect 2177 632 2518 678
rect 2177 590 2223 632
rect 1834 308 1907 354
rect 1834 262 1845 308
rect 1891 262 1907 308
rect 1834 261 1907 262
rect 2177 215 2223 544
rect 1742 169 1933 215
rect 1979 169 1990 215
rect 1573 158 1696 169
rect 2177 156 2223 169
rect 2269 574 2415 585
rect 2269 528 2369 574
rect 2269 515 2415 528
rect 2472 523 2518 632
rect 2581 615 2650 724
rect 2581 569 2593 615
rect 2639 569 2650 615
rect 2700 632 3067 678
rect 2700 523 2746 632
rect 2269 348 2319 515
rect 2472 476 2746 523
rect 2797 574 2843 585
rect 2367 414 2747 426
rect 2367 368 2682 414
rect 2728 368 2747 414
rect 2367 356 2747 368
rect 2269 302 2270 348
rect 2316 302 2319 348
rect 2269 229 2319 302
rect 2269 216 2415 229
rect 2269 170 2349 216
rect 2395 170 2415 216
rect 2269 159 2415 170
rect 2573 216 2619 229
rect 2573 60 2619 170
rect 2797 216 2843 528
rect 2797 156 2843 170
rect 3001 574 3067 632
rect 3438 609 3506 724
rect 3047 528 3067 574
rect 3001 216 3067 528
rect 3001 170 3021 216
rect 3113 563 3228 609
rect 3274 563 3285 609
rect 3438 563 3449 609
rect 3495 563 3506 609
rect 3672 609 3739 628
rect 3672 563 3673 609
rect 3719 563 3739 609
rect 3113 216 3159 563
rect 3672 517 3739 563
rect 3205 471 3739 517
rect 3205 392 3251 471
rect 3297 412 3635 424
rect 3297 366 3353 412
rect 3399 366 3635 412
rect 3297 356 3635 366
rect 3205 335 3251 346
rect 3469 216 3515 229
rect 3113 170 3245 216
rect 3291 170 3302 216
rect 3001 156 3067 170
rect 3469 60 3515 170
rect 3693 216 3739 471
rect 3693 156 3739 170
rect 0 -60 3808 60
<< labels >>
flabel metal1 s 3297 356 3635 424 0 FreeSans 400 0 0 0 I0
port 1 nsew default input
flabel metal1 s 1481 229 1527 232 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 0 724 3808 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 141 194 202 590 0 FreeSans 400 0 0 0 I2
port 3 nsew default input
flabel metal1 s 2367 356 2747 426 0 FreeSans 400 0 0 0 I1
port 2 nsew default input
flabel metal1 s 451 360 740 450 0 FreeSans 400 0 0 0 S0
port 5 nsew default input
flabel metal1 s 901 360 1151 430 0 FreeSans 400 0 0 0 I3
port 4 nsew default input
flabel metal1 s 2033 430 2107 664 0 FreeSans 400 0 0 0 S1
port 6 nsew default input
flabel metal1 s 1246 120 1320 571 0 FreeSans 400 0 0 0 Z
port 7 nsew default output
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 901 110 987 360 1 I3
port 4 nsew default input
rlabel metal1 s 660 248 740 360 1 S0
port 5 nsew default input
rlabel metal1 s 1834 354 2107 430 1 S1
port 6 nsew default input
rlabel metal1 s 1834 261 1907 354 1 S1
port 6 nsew default input
rlabel metal1 s 3438 569 3506 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2581 569 2650 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1481 569 1527 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1002 569 1070 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 569 95 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3438 563 3506 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1481 563 1527 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 563 95 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1481 515 1527 563 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 49 515 95 563 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1481 514 1527 515 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1033 229 1079 232 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3469 226 3515 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2573 226 2619 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1481 226 1527 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1033 226 1079 229 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 3469 60 3515 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2573 60 2619 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1481 60 1527 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1033 60 1079 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 226 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string GDS_END 677056
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 669126
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
