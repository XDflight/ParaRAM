magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -64 2204 65 2243
rect -64 2148 -28 2204
rect 28 2148 65 2204
rect -64 1987 65 2148
rect -64 1931 -28 1987
rect 28 1931 65 1987
rect -64 1769 65 1931
rect -64 1713 -28 1769
rect 28 1713 65 1769
rect -64 1551 65 1713
rect -64 1495 -28 1551
rect 28 1495 65 1551
rect -64 1334 65 1495
rect -64 1278 -28 1334
rect 28 1278 65 1334
rect -64 1116 65 1278
rect -64 1060 -28 1116
rect 28 1060 65 1116
rect -64 899 65 1060
rect -64 843 -28 899
rect 28 843 65 899
rect -64 681 65 843
rect -64 625 -28 681
rect 28 625 65 681
rect -64 463 65 625
rect -64 407 -28 463
rect 28 407 65 463
rect -64 246 65 407
rect -64 190 -28 246
rect 28 190 65 246
rect -64 28 65 190
rect -64 -28 -28 28
rect 28 -28 65 28
rect -64 -190 65 -28
rect -64 -246 -28 -190
rect 28 -246 65 -190
rect -64 -407 65 -246
rect -64 -463 -28 -407
rect 28 -463 65 -407
rect -64 -625 65 -463
rect -64 -681 -28 -625
rect 28 -681 65 -625
rect -64 -843 65 -681
rect -64 -899 -28 -843
rect 28 -899 65 -843
rect -64 -1060 65 -899
rect -64 -1116 -28 -1060
rect 28 -1116 65 -1060
rect -64 -1278 65 -1116
rect -64 -1334 -28 -1278
rect 28 -1334 65 -1278
rect -64 -1495 65 -1334
rect -64 -1551 -28 -1495
rect 28 -1551 65 -1495
rect -64 -1713 65 -1551
rect -64 -1769 -28 -1713
rect 28 -1769 65 -1713
rect -64 -1931 65 -1769
rect -64 -1987 -28 -1931
rect 28 -1987 65 -1931
rect -64 -2148 65 -1987
rect -64 -2204 -28 -2148
rect 28 -2204 65 -2148
rect -64 -2243 65 -2204
<< via2 >>
rect -28 2148 28 2204
rect -28 1931 28 1987
rect -28 1713 28 1769
rect -28 1495 28 1551
rect -28 1278 28 1334
rect -28 1060 28 1116
rect -28 843 28 899
rect -28 625 28 681
rect -28 407 28 463
rect -28 190 28 246
rect -28 -28 28 28
rect -28 -246 28 -190
rect -28 -463 28 -407
rect -28 -681 28 -625
rect -28 -899 28 -843
rect -28 -1116 28 -1060
rect -28 -1334 28 -1278
rect -28 -1551 28 -1495
rect -28 -1769 28 -1713
rect -28 -1987 28 -1931
rect -28 -2204 28 -2148
<< metal3 >>
rect -65 2204 65 2243
rect -65 2148 -28 2204
rect 28 2148 65 2204
rect -65 1987 65 2148
rect -65 1931 -28 1987
rect 28 1931 65 1987
rect -65 1769 65 1931
rect -65 1713 -28 1769
rect 28 1713 65 1769
rect -65 1551 65 1713
rect -65 1495 -28 1551
rect 28 1495 65 1551
rect -65 1334 65 1495
rect -65 1278 -28 1334
rect 28 1278 65 1334
rect -65 1116 65 1278
rect -65 1060 -28 1116
rect 28 1060 65 1116
rect -65 899 65 1060
rect -65 843 -28 899
rect 28 843 65 899
rect -65 681 65 843
rect -65 625 -28 681
rect 28 625 65 681
rect -65 463 65 625
rect -65 407 -28 463
rect 28 407 65 463
rect -65 246 65 407
rect -65 190 -28 246
rect 28 190 65 246
rect -65 28 65 190
rect -65 -28 -28 28
rect 28 -28 65 28
rect -65 -190 65 -28
rect -65 -246 -28 -190
rect 28 -246 65 -190
rect -65 -407 65 -246
rect -65 -463 -28 -407
rect 28 -463 65 -407
rect -65 -625 65 -463
rect -65 -681 -28 -625
rect 28 -681 65 -625
rect -65 -843 65 -681
rect -65 -899 -28 -843
rect 28 -899 65 -843
rect -65 -1060 65 -899
rect -65 -1116 -28 -1060
rect 28 -1116 65 -1060
rect -65 -1278 65 -1116
rect -65 -1334 -28 -1278
rect 28 -1334 65 -1278
rect -65 -1495 65 -1334
rect -65 -1551 -28 -1495
rect 28 -1551 65 -1495
rect -65 -1713 65 -1551
rect -65 -1769 -28 -1713
rect 28 -1769 65 -1713
rect -65 -1931 65 -1769
rect -65 -1987 -28 -1931
rect 28 -1987 65 -1931
rect -65 -2148 65 -1987
rect -65 -2204 -28 -2148
rect 28 -2204 65 -2148
rect -65 -2243 65 -2204
<< properties >>
string GDS_END 1106730
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1105254
<< end >>
