magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 682
rect 224 0 344 682
rect 448 0 568 682
rect 672 0 792 682
rect 896 0 1016 682
rect 1120 0 1240 682
rect 1344 0 1464 682
rect 1568 0 1688 682
<< mvndiff >>
rect -88 669 0 682
rect -88 13 -75 669
rect -29 13 0 669
rect -88 0 0 13
rect 120 669 224 682
rect 120 13 149 669
rect 195 13 224 669
rect 120 0 224 13
rect 344 669 448 682
rect 344 13 373 669
rect 419 13 448 669
rect 344 0 448 13
rect 568 669 672 682
rect 568 13 597 669
rect 643 13 672 669
rect 568 0 672 13
rect 792 669 896 682
rect 792 13 821 669
rect 867 13 896 669
rect 792 0 896 13
rect 1016 669 1120 682
rect 1016 13 1045 669
rect 1091 13 1120 669
rect 1016 0 1120 13
rect 1240 669 1344 682
rect 1240 13 1269 669
rect 1315 13 1344 669
rect 1240 0 1344 13
rect 1464 669 1568 682
rect 1464 13 1493 669
rect 1539 13 1568 669
rect 1464 0 1568 13
rect 1688 669 1776 682
rect 1688 13 1717 669
rect 1763 13 1776 669
rect 1688 0 1776 13
<< mvndiffc >>
rect -75 13 -29 669
rect 149 13 195 669
rect 373 13 419 669
rect 597 13 643 669
rect 821 13 867 669
rect 1045 13 1091 669
rect 1269 13 1315 669
rect 1493 13 1539 669
rect 1717 13 1763 669
<< polysilicon >>
rect 0 682 120 726
rect 224 682 344 726
rect 448 682 568 726
rect 672 682 792 726
rect 896 682 1016 726
rect 1120 682 1240 726
rect 1344 682 1464 726
rect 1568 682 1688 726
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
<< metal1 >>
rect -75 669 -29 682
rect -75 0 -29 13
rect 149 669 195 682
rect 149 0 195 13
rect 373 669 419 682
rect 373 0 419 13
rect 597 669 643 682
rect 597 0 643 13
rect 821 669 867 682
rect 821 0 867 13
rect 1045 669 1091 682
rect 1045 0 1091 13
rect 1269 669 1315 682
rect 1269 0 1315 13
rect 1493 669 1539 682
rect 1493 0 1539 13
rect 1717 669 1763 682
rect 1717 0 1763 13
<< labels >>
flabel metal1 s -52 341 -52 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 1740 341 1740 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 341 172 341 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 341 396 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 341 620 341 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 341 844 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 341 1068 341 0 FreeSans 200 0 0 0 D
flabel metal1 s 1292 341 1292 341 0 FreeSans 200 0 0 0 S
flabel metal1 s 1516 341 1516 341 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 64174
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 56572
<< end >>
