magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -50 169 50 174
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -174 50 -169
<< via2 >>
rect -45 141 -17 169
rect 17 141 45 169
rect -45 79 -17 107
rect 17 79 45 107
rect -45 17 -17 45
rect 17 17 45 45
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect -45 -169 -17 -141
rect 17 -169 45 -141
<< metal3 >>
rect -50 169 50 174
rect -50 141 -45 169
rect -17 141 17 169
rect 45 141 50 169
rect -50 107 50 141
rect -50 79 -45 107
rect -17 79 17 107
rect 45 79 50 107
rect -50 45 50 79
rect -50 17 -45 45
rect -17 17 17 45
rect 45 17 50 45
rect -50 -17 50 17
rect -50 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 50 -17
rect -50 -79 50 -45
rect -50 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 50 -79
rect -50 -141 50 -107
rect -50 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 50 -141
rect -50 -174 50 -169
<< properties >>
string GDS_END 664600
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 663700
<< end >>
