magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 328 3658
<< mvpmos >>
rect 0 0 120 3538
<< mvpdiff >>
rect -88 3525 0 3538
rect -88 13 -75 3525
rect -29 13 0 3525
rect -88 0 0 13
rect 120 3525 208 3538
rect 120 13 149 3525
rect 195 13 208 3525
rect 120 0 208 13
<< mvpdiffc >>
rect -75 13 -29 3525
rect 149 13 195 3525
<< polysilicon >>
rect 0 3538 120 3582
rect 0 -44 120 0
<< metal1 >>
rect -75 3525 -29 3538
rect -75 0 -29 13
rect 149 3525 195 3538
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1769 -52 1769 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1769 172 1769 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 113840
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 108400
<< end >>
