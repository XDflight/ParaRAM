magic
tech gf180mcuA
timestamp 1666464484
<< metal1 >>
rect 0 147 78 159
rect 13 106 18 147
rect 42 99 47 140
rect 59 106 64 147
rect 42 93 67 99
rect 29 80 39 86
rect 9 67 19 73
rect 44 67 54 73
rect 59 47 64 93
rect 59 42 66 47
rect 27 9 32 27
rect 61 16 66 42
rect 0 -3 78 9
<< obsm1 >>
rect 10 32 49 37
rect 10 16 15 32
rect 44 16 49 32
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 9 148 19 154
rect 33 148 43 154
rect 57 148 67 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 57 92 67 100
rect 29 79 39 87
rect 9 66 19 74
rect 44 66 54 74
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 9 2 19 8
rect 33 2 43 8
rect 57 2 67 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
<< labels >>
rlabel metal2 s 9 66 19 74 6 A0
port 1 nsew signal input
rlabel metal1 s 9 67 19 73 6 A0
port 1 nsew signal input
rlabel metal2 s 29 79 39 87 6 A1
port 2 nsew signal input
rlabel metal1 s 29 80 39 86 6 A1
port 2 nsew signal input
rlabel metal2 s 44 66 54 74 6 B
port 3 nsew signal input
rlabel metal1 s 44 67 54 73 6 B
port 3 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 34 147 42 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 33 148 43 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 58 147 66 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 57 148 67 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 13 106 18 159 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 59 106 64 159 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 147 78 159 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 34 1 42 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 33 2 43 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 58 1 66 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 57 2 67 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 27 -3 32 27 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 0 -3 78 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 57 92 67 100 6 Y
port 6 nsew signal output
rlabel metal1 s 42 93 47 140 6 Y
port 6 nsew signal output
rlabel metal1 s 59 42 64 99 6 Y
port 6 nsew signal output
rlabel metal1 s 61 16 66 47 6 Y
port 6 nsew signal output
rlabel metal1 s 42 93 67 99 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 78 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
