magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -2204 23 2204 42
rect -2204 -23 -2185 23
rect 2185 -23 2204 23
rect -2204 -42 2204 -23
<< polycontact >>
rect -2185 -23 2185 23
<< metal1 >>
rect -2196 23 2196 34
rect -2196 -23 -2185 23
rect 2185 -23 2196 23
rect -2196 -34 2196 -23
<< properties >>
string GDS_END 1004888
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1001748
<< end >>
