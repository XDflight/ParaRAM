magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1430 1094
<< pwell >>
rect -86 -86 1430 453
<< mvnmos >>
rect 124 69 244 279
rect 348 69 468 279
rect 572 69 692 279
rect 832 69 952 333
rect 1056 69 1176 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 842 573 942 939
rect 1056 573 1156 939
<< mvndiff >>
rect 752 279 832 333
rect 36 193 124 279
rect 36 147 49 193
rect 95 147 124 193
rect 36 69 124 147
rect 244 266 348 279
rect 244 126 273 266
rect 319 126 348 266
rect 244 69 348 126
rect 468 193 572 279
rect 468 147 497 193
rect 543 147 572 193
rect 468 69 572 147
rect 692 266 832 279
rect 692 126 721 266
rect 767 126 832 266
rect 692 69 832 126
rect 952 287 1056 333
rect 952 147 981 287
rect 1027 147 1056 287
rect 952 69 1056 147
rect 1176 287 1264 333
rect 1176 147 1205 287
rect 1251 147 1264 287
rect 1176 69 1264 147
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 573 582 939
rect 682 861 842 939
rect 682 721 711 861
rect 757 721 842 861
rect 682 573 842 721
rect 942 861 1056 939
rect 942 721 971 861
rect 1017 721 1056 861
rect 942 573 1056 721
rect 1156 861 1244 939
rect 1156 721 1185 861
rect 1231 721 1244 861
rect 1156 573 1244 721
<< mvndiffc >>
rect 49 147 95 193
rect 273 126 319 266
rect 497 147 543 193
rect 721 126 767 266
rect 981 147 1027 287
rect 1205 147 1251 287
<< mvpdiffc >>
rect 69 721 115 861
rect 711 721 757 861
rect 971 721 1017 861
rect 1185 721 1231 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 842 939 942 983
rect 1056 939 1156 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 323 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 323 458 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 323 682 454
rect 842 513 942 573
rect 1056 513 1156 573
rect 842 500 1156 513
rect 842 454 855 500
rect 901 454 1156 500
rect 842 441 1156 454
rect 842 377 952 441
rect 832 333 952 377
rect 1056 377 1156 441
rect 1056 333 1176 377
rect 124 279 244 323
rect 348 279 468 323
rect 572 279 692 323
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 832 25 952 69
rect 1056 25 1176 69
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 595 454 641 500
rect 855 454 901 500
<< metal1 >>
rect 0 918 1344 1098
rect 69 861 115 872
rect 69 664 115 721
rect 711 861 757 918
rect 711 710 757 721
rect 926 861 1027 872
rect 926 721 971 861
rect 1017 721 1027 861
rect 69 618 734 664
rect 142 500 214 542
rect 142 454 157 500
rect 203 454 214 500
rect 359 500 418 542
rect 359 454 371 500
rect 417 454 418 500
rect 359 443 418 454
rect 583 500 642 542
rect 583 454 595 500
rect 641 454 642 500
rect 583 443 642 454
rect 688 511 734 618
rect 926 578 1027 721
rect 1185 861 1231 918
rect 1185 710 1231 721
rect 688 500 901 511
rect 688 454 855 500
rect 688 443 901 454
rect 688 369 734 443
rect 49 323 734 369
rect 49 193 95 323
rect 49 136 95 147
rect 273 266 319 277
rect 497 193 543 323
rect 981 287 1027 578
rect 497 136 543 147
rect 721 266 767 277
rect 273 90 319 126
rect 981 136 1027 147
rect 1205 287 1251 298
rect 721 90 767 126
rect 1205 90 1251 147
rect 0 -90 1344 90
<< labels >>
flabel metal1 s 142 454 214 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 359 443 418 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 583 443 642 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 918 1344 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1205 277 1251 298 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 926 578 1027 872 0 FreeSans 200 0 0 0 Z
port 4 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 981 136 1027 578 1 Z
port 4 nsew default output
rlabel metal1 s 1185 710 1231 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 711 710 757 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1205 90 1251 277 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 721 90 767 277 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 277 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1344 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 1008
string GDS_END 276230
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 272340
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
