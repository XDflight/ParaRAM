magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 328 3160
<< mvpmos >>
rect 0 0 120 3040
<< mvpdiff >>
rect -88 3027 0 3040
rect -88 1043 -75 3027
rect -29 1043 0 3027
rect -88 986 0 1043
rect -88 940 -75 986
rect -29 940 0 986
rect -88 883 0 940
rect -88 837 -75 883
rect -29 837 0 883
rect -88 780 0 837
rect -88 734 -75 780
rect -29 734 0 780
rect -88 677 0 734
rect -88 631 -75 677
rect -29 631 0 677
rect -88 574 0 631
rect -88 528 -75 574
rect -29 528 0 574
rect -88 471 0 528
rect -88 425 -75 471
rect -29 425 0 471
rect -88 368 0 425
rect -88 322 -75 368
rect -29 322 0 368
rect -88 265 0 322
rect -88 219 -75 265
rect -29 219 0 265
rect -88 162 0 219
rect -88 116 -75 162
rect -29 116 0 162
rect -88 59 0 116
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 3027 208 3040
rect 120 1043 149 3027
rect 195 1043 208 3027
rect 120 986 208 1043
rect 120 940 149 986
rect 195 940 208 986
rect 120 883 208 940
rect 120 837 149 883
rect 195 837 208 883
rect 120 780 208 837
rect 120 734 149 780
rect 195 734 208 780
rect 120 677 208 734
rect 120 631 149 677
rect 195 631 208 677
rect 120 574 208 631
rect 120 528 149 574
rect 195 528 208 574
rect 120 471 208 528
rect 120 425 149 471
rect 195 425 208 471
rect 120 368 208 425
rect 120 322 149 368
rect 195 322 208 368
rect 120 265 208 322
rect 120 219 149 265
rect 195 219 208 265
rect 120 162 208 219
rect 120 116 149 162
rect 195 116 208 162
rect 120 59 208 116
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvpdiffc >>
rect -75 1043 -29 3027
rect -75 940 -29 986
rect -75 837 -29 883
rect -75 734 -29 780
rect -75 631 -29 677
rect -75 528 -29 574
rect -75 425 -29 471
rect -75 322 -29 368
rect -75 219 -29 265
rect -75 116 -29 162
rect -75 13 -29 59
rect 149 1043 195 3027
rect 149 940 195 986
rect 149 837 195 883
rect 149 734 195 780
rect 149 631 195 677
rect 149 528 195 574
rect 149 425 195 471
rect 149 322 195 368
rect 149 219 195 265
rect 149 116 195 162
rect 149 13 195 59
<< polysilicon >>
rect 0 3040 120 3084
rect 0 -44 120 0
<< metal1 >>
rect -75 3027 -29 3040
rect -75 986 -29 1043
rect -75 883 -29 940
rect -75 780 -29 837
rect -75 677 -29 734
rect -75 574 -29 631
rect -75 471 -29 528
rect -75 368 -29 425
rect -75 265 -29 322
rect -75 162 -29 219
rect -75 59 -29 116
rect -75 0 -29 13
rect 149 3027 195 3040
rect 149 986 195 1043
rect 149 883 195 940
rect 149 780 195 837
rect 149 677 195 734
rect 149 574 195 631
rect 149 471 195 528
rect 149 368 195 425
rect 149 265 195 322
rect 149 162 195 219
rect 149 59 195 116
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 1520 -52 1520 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1520 172 1520 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 41062
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 36262
<< end >>
