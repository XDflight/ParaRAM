magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 874
<< mvpmos >>
rect 0 0 120 754
rect 224 0 344 754
<< mvpdiff >>
rect -88 741 0 754
rect -88 695 -75 741
rect -29 695 0 741
rect -88 628 0 695
rect -88 582 -75 628
rect -29 582 0 628
rect -88 515 0 582
rect -88 469 -75 515
rect -29 469 0 515
rect -88 401 0 469
rect -88 355 -75 401
rect -29 355 0 401
rect -88 287 0 355
rect -88 241 -75 287
rect -29 241 0 287
rect -88 173 0 241
rect -88 127 -75 173
rect -29 127 0 173
rect -88 59 0 127
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 741 224 754
rect 120 695 149 741
rect 195 695 224 741
rect 120 628 224 695
rect 120 582 149 628
rect 195 582 224 628
rect 120 515 224 582
rect 120 469 149 515
rect 195 469 224 515
rect 120 401 224 469
rect 120 355 149 401
rect 195 355 224 401
rect 120 287 224 355
rect 120 241 149 287
rect 195 241 224 287
rect 120 173 224 241
rect 120 127 149 173
rect 195 127 224 173
rect 120 59 224 127
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 741 432 754
rect 344 695 373 741
rect 419 695 432 741
rect 344 628 432 695
rect 344 582 373 628
rect 419 582 432 628
rect 344 515 432 582
rect 344 469 373 515
rect 419 469 432 515
rect 344 401 432 469
rect 344 355 373 401
rect 419 355 432 401
rect 344 287 432 355
rect 344 241 373 287
rect 419 241 432 287
rect 344 173 432 241
rect 344 127 373 173
rect 419 127 432 173
rect 344 59 432 127
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 695 -29 741
rect -75 582 -29 628
rect -75 469 -29 515
rect -75 355 -29 401
rect -75 241 -29 287
rect -75 127 -29 173
rect -75 13 -29 59
rect 149 695 195 741
rect 149 582 195 628
rect 149 469 195 515
rect 149 355 195 401
rect 149 241 195 287
rect 149 127 195 173
rect 149 13 195 59
rect 373 695 419 741
rect 373 582 419 628
rect 373 469 419 515
rect 373 355 419 401
rect 373 241 419 287
rect 373 127 419 173
rect 373 13 419 59
<< polysilicon >>
rect 0 754 120 798
rect 224 754 344 798
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 741 -29 754
rect -75 628 -29 695
rect -75 515 -29 582
rect -75 401 -29 469
rect -75 287 -29 355
rect -75 173 -29 241
rect -75 59 -29 127
rect -75 0 -29 13
rect 149 741 195 754
rect 149 628 195 695
rect 149 515 195 582
rect 149 401 195 469
rect 149 287 195 355
rect 149 173 195 241
rect 149 59 195 127
rect 149 0 195 13
rect 373 741 419 754
rect 373 628 419 695
rect 373 515 419 582
rect 373 401 419 469
rect 373 287 419 355
rect 373 173 419 241
rect 373 59 419 127
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 377 -52 377 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 377 396 377 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 377 172 377 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 523768
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 521082
<< end >>
