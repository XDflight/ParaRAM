magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 1448 876
<< mvpmos >>
rect 0 0 120 756
rect 224 0 344 756
rect 448 0 568 756
rect 672 0 792 756
rect 896 0 1016 756
rect 1120 0 1240 756
<< mvpdiff >>
rect -88 743 0 756
rect -88 697 -75 743
rect -29 697 0 743
rect -88 629 0 697
rect -88 583 -75 629
rect -29 583 0 629
rect -88 515 0 583
rect -88 469 -75 515
rect -29 469 0 515
rect -88 401 0 469
rect -88 355 -75 401
rect -29 355 0 401
rect -88 287 0 355
rect -88 241 -75 287
rect -29 241 0 287
rect -88 173 0 241
rect -88 127 -75 173
rect -29 127 0 173
rect -88 59 0 127
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 743 224 756
rect 120 697 149 743
rect 195 697 224 743
rect 120 629 224 697
rect 120 583 149 629
rect 195 583 224 629
rect 120 515 224 583
rect 120 469 149 515
rect 195 469 224 515
rect 120 401 224 469
rect 120 355 149 401
rect 195 355 224 401
rect 120 287 224 355
rect 120 241 149 287
rect 195 241 224 287
rect 120 173 224 241
rect 120 127 149 173
rect 195 127 224 173
rect 120 59 224 127
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 743 448 756
rect 344 697 373 743
rect 419 697 448 743
rect 344 629 448 697
rect 344 583 373 629
rect 419 583 448 629
rect 344 515 448 583
rect 344 469 373 515
rect 419 469 448 515
rect 344 401 448 469
rect 344 355 373 401
rect 419 355 448 401
rect 344 287 448 355
rect 344 241 373 287
rect 419 241 448 287
rect 344 173 448 241
rect 344 127 373 173
rect 419 127 448 173
rect 344 59 448 127
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 743 672 756
rect 568 697 597 743
rect 643 697 672 743
rect 568 629 672 697
rect 568 583 597 629
rect 643 583 672 629
rect 568 515 672 583
rect 568 469 597 515
rect 643 469 672 515
rect 568 401 672 469
rect 568 355 597 401
rect 643 355 672 401
rect 568 287 672 355
rect 568 241 597 287
rect 643 241 672 287
rect 568 173 672 241
rect 568 127 597 173
rect 643 127 672 173
rect 568 59 672 127
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 743 896 756
rect 792 697 821 743
rect 867 697 896 743
rect 792 629 896 697
rect 792 583 821 629
rect 867 583 896 629
rect 792 515 896 583
rect 792 469 821 515
rect 867 469 896 515
rect 792 401 896 469
rect 792 355 821 401
rect 867 355 896 401
rect 792 287 896 355
rect 792 241 821 287
rect 867 241 896 287
rect 792 173 896 241
rect 792 127 821 173
rect 867 127 896 173
rect 792 59 896 127
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 743 1120 756
rect 1016 697 1045 743
rect 1091 697 1120 743
rect 1016 629 1120 697
rect 1016 583 1045 629
rect 1091 583 1120 629
rect 1016 515 1120 583
rect 1016 469 1045 515
rect 1091 469 1120 515
rect 1016 401 1120 469
rect 1016 355 1045 401
rect 1091 355 1120 401
rect 1016 287 1120 355
rect 1016 241 1045 287
rect 1091 241 1120 287
rect 1016 173 1120 241
rect 1016 127 1045 173
rect 1091 127 1120 173
rect 1016 59 1120 127
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 743 1328 756
rect 1240 697 1269 743
rect 1315 697 1328 743
rect 1240 629 1328 697
rect 1240 583 1269 629
rect 1315 583 1328 629
rect 1240 515 1328 583
rect 1240 469 1269 515
rect 1315 469 1328 515
rect 1240 401 1328 469
rect 1240 355 1269 401
rect 1315 355 1328 401
rect 1240 287 1328 355
rect 1240 241 1269 287
rect 1315 241 1328 287
rect 1240 173 1328 241
rect 1240 127 1269 173
rect 1315 127 1328 173
rect 1240 59 1328 127
rect 1240 13 1269 59
rect 1315 13 1328 59
rect 1240 0 1328 13
<< mvpdiffc >>
rect -75 697 -29 743
rect -75 583 -29 629
rect -75 469 -29 515
rect -75 355 -29 401
rect -75 241 -29 287
rect -75 127 -29 173
rect -75 13 -29 59
rect 149 697 195 743
rect 149 583 195 629
rect 149 469 195 515
rect 149 355 195 401
rect 149 241 195 287
rect 149 127 195 173
rect 149 13 195 59
rect 373 697 419 743
rect 373 583 419 629
rect 373 469 419 515
rect 373 355 419 401
rect 373 241 419 287
rect 373 127 419 173
rect 373 13 419 59
rect 597 697 643 743
rect 597 583 643 629
rect 597 469 643 515
rect 597 355 643 401
rect 597 241 643 287
rect 597 127 643 173
rect 597 13 643 59
rect 821 697 867 743
rect 821 583 867 629
rect 821 469 867 515
rect 821 355 867 401
rect 821 241 867 287
rect 821 127 867 173
rect 821 13 867 59
rect 1045 697 1091 743
rect 1045 583 1091 629
rect 1045 469 1091 515
rect 1045 355 1091 401
rect 1045 241 1091 287
rect 1045 127 1091 173
rect 1045 13 1091 59
rect 1269 697 1315 743
rect 1269 583 1315 629
rect 1269 469 1315 515
rect 1269 355 1315 401
rect 1269 241 1315 287
rect 1269 127 1315 173
rect 1269 13 1315 59
<< polysilicon >>
rect 0 756 120 800
rect 224 756 344 800
rect 448 756 568 800
rect 672 756 792 800
rect 896 756 1016 800
rect 1120 756 1240 800
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
<< metal1 >>
rect -75 743 -29 756
rect -75 629 -29 697
rect -75 515 -29 583
rect -75 401 -29 469
rect -75 287 -29 355
rect -75 173 -29 241
rect -75 59 -29 127
rect -75 0 -29 13
rect 149 743 195 756
rect 149 629 195 697
rect 149 515 195 583
rect 149 401 195 469
rect 149 287 195 355
rect 149 173 195 241
rect 149 59 195 127
rect 149 0 195 13
rect 373 743 419 756
rect 373 629 419 697
rect 373 515 419 583
rect 373 401 419 469
rect 373 287 419 355
rect 373 173 419 241
rect 373 59 419 127
rect 373 0 419 13
rect 597 743 643 756
rect 597 629 643 697
rect 597 515 643 583
rect 597 401 643 469
rect 597 287 643 355
rect 597 173 643 241
rect 597 59 643 127
rect 597 0 643 13
rect 821 743 867 756
rect 821 629 867 697
rect 821 515 867 583
rect 821 401 867 469
rect 821 287 867 355
rect 821 173 867 241
rect 821 59 867 127
rect 821 0 867 13
rect 1045 743 1091 756
rect 1045 629 1091 697
rect 1045 515 1091 583
rect 1045 401 1091 469
rect 1045 287 1091 355
rect 1045 173 1091 241
rect 1045 59 1091 127
rect 1045 0 1091 13
rect 1269 743 1315 756
rect 1269 629 1315 697
rect 1269 515 1315 583
rect 1269 401 1315 469
rect 1269 287 1315 355
rect 1269 173 1315 241
rect 1269 59 1315 127
rect 1269 0 1315 13
<< labels >>
flabel metal1 s -52 378 -52 378 0 FreeSans 400 0 0 0 S
flabel metal1 s 1292 378 1292 378 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 378 172 378 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 378 396 378 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 378 620 378 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 378 844 378 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 378 1068 378 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 225268
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 219262
<< end >>
