magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -203 10266 787 12370
rect -7 8752 622 10266
rect -7 8695 624 8752
rect -5 7108 624 8695
rect -221 1164 756 1620
rect -203 648 756 1164
<< pmos >>
rect 138 11191 258 11873
rect 362 11191 482 11873
rect 138 10416 258 11098
rect 362 10416 482 11098
rect 67 788 187 1085
rect 319 788 439 1085
<< pdiff >>
rect 0 11828 138 11873
rect 23 11782 138 11828
rect 0 11646 138 11782
rect 23 11600 138 11646
rect 0 11465 138 11600
rect 23 11419 138 11465
rect 0 11283 138 11419
rect 23 11237 138 11283
rect 0 11191 138 11237
rect 258 11828 362 11873
rect 258 11782 287 11828
rect 333 11782 362 11828
rect 258 11646 362 11782
rect 258 11600 287 11646
rect 333 11600 362 11646
rect 258 11465 362 11600
rect 258 11419 287 11465
rect 333 11419 362 11465
rect 258 11283 362 11419
rect 258 11237 287 11283
rect 333 11237 362 11283
rect 258 11191 362 11237
rect 482 11828 650 11873
rect 482 11782 513 11828
rect 559 11782 650 11828
rect 482 11646 650 11782
rect 482 11600 513 11646
rect 559 11600 650 11646
rect 482 11465 650 11600
rect 482 11419 513 11465
rect 559 11419 650 11465
rect 482 11283 650 11419
rect 482 11237 513 11283
rect 559 11237 650 11283
rect 482 11191 650 11237
rect 0 11052 138 11098
rect 23 11006 138 11052
rect 0 10871 138 11006
rect 23 10825 138 10871
rect 0 10690 138 10825
rect 23 10644 138 10690
rect 0 10508 138 10644
rect 23 10462 138 10508
rect 0 10416 138 10462
rect 258 11052 362 11098
rect 258 11006 287 11052
rect 333 11006 362 11052
rect 258 10871 362 11006
rect 258 10825 287 10871
rect 333 10825 362 10871
rect 258 10690 362 10825
rect 258 10644 287 10690
rect 333 10644 362 10690
rect 258 10508 362 10644
rect 258 10462 287 10508
rect 333 10462 362 10508
rect 258 10416 362 10462
rect 482 11052 650 11098
rect 482 11006 513 11052
rect 559 11006 650 11052
rect 482 10871 650 11006
rect 482 10825 513 10871
rect 559 10825 650 10871
rect 482 10690 650 10825
rect 482 10644 513 10690
rect 559 10644 650 10690
rect 482 10508 650 10644
rect 482 10462 513 10508
rect 559 10462 650 10508
rect 482 10416 650 10462
rect -67 960 67 1085
rect -67 914 -23 960
rect 23 914 67 960
rect -67 788 67 914
rect 187 960 319 1085
rect 187 914 230 960
rect 276 914 319 960
rect 187 788 319 914
rect 439 960 620 1085
rect 439 914 480 960
rect 526 914 620 960
rect 439 788 620 914
<< pdiffc >>
rect -1 11782 23 11828
rect -1 11600 23 11646
rect -1 11419 23 11465
rect -1 11237 23 11283
rect 287 11782 333 11828
rect 287 11600 333 11646
rect 287 11419 333 11465
rect 287 11237 333 11283
rect 513 11782 559 11828
rect 513 11600 559 11646
rect 513 11419 559 11465
rect 513 11237 559 11283
rect -1 11006 23 11052
rect -1 10825 23 10871
rect -1 10644 23 10690
rect -1 10462 23 10508
rect 287 11006 333 11052
rect 287 10825 333 10871
rect 287 10644 333 10690
rect 287 10462 333 10508
rect 513 11006 559 11052
rect 513 10825 559 10871
rect 513 10644 559 10690
rect 513 10462 559 10508
rect -23 914 23 960
rect 230 914 276 960
rect 480 914 526 960
<< psubdiff >>
rect -80 5260 80 5320
rect -80 5214 -23 5260
rect 23 5214 80 5260
rect -80 5154 80 5214
rect -80 96 620 155
rect -80 50 -23 96
rect 23 50 135 96
rect 181 50 293 96
rect 339 50 451 96
rect 497 50 620 96
rect -80 -10 620 50
<< nsubdiff >>
rect -1 12165 650 12222
rect -1 12119 129 12165
rect 175 12119 287 12165
rect 333 12119 445 12165
rect 491 12119 650 12165
rect -1 12062 650 12119
rect -78 1415 620 1472
rect -78 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -78 1312 620 1369
<< psubdiffcont >>
rect -23 5214 23 5260
rect -23 50 23 96
rect 135 50 181 96
rect 293 50 339 96
rect 451 50 497 96
<< nsubdiffcont >>
rect 129 12119 175 12165
rect 287 12119 333 12165
rect 445 12119 491 12165
rect -23 1369 23 1415
rect 135 1369 181 1415
rect 293 1369 339 1415
rect 451 1369 497 1415
<< polysilicon >>
rect 138 11873 258 11946
rect 362 11873 482 11946
rect 138 11098 258 11191
rect 362 11098 482 11191
rect 138 10352 258 10416
rect 362 10352 482 10416
rect 138 10333 482 10352
rect 138 10287 170 10333
rect 404 10287 482 10333
rect 138 10268 482 10287
rect 248 10198 368 10268
rect 248 8764 368 8836
rect 250 8611 370 8684
rect 250 7164 370 7249
rect 250 7118 293 7164
rect 339 7118 370 7164
rect 250 7099 370 7118
rect 250 4968 369 5505
rect 250 3469 370 3516
rect 250 3423 287 3469
rect 333 3423 370 3469
rect 250 3404 370 3423
rect 250 3192 370 3211
rect 250 3146 287 3192
rect 333 3146 370 3192
rect 250 3099 370 3146
rect 67 1225 439 1244
rect 67 1179 230 1225
rect 276 1179 439 1225
rect 67 1145 439 1179
rect 67 1085 187 1145
rect 319 1085 439 1145
rect 67 661 187 788
rect 67 612 172 661
rect 52 539 172 612
rect 319 601 439 788
rect 319 570 396 601
rect 276 539 396 570
rect 52 497 170 498
rect 52 310 172 382
rect 276 310 396 382
<< polycontact >>
rect 170 10287 404 10333
rect 293 7118 339 7164
rect 287 3423 333 3469
rect 287 3146 333 3192
rect 230 1179 276 1225
<< metal1 >>
rect -58 12203 620 12227
rect -58 12165 281 12203
rect 333 12165 620 12203
rect -58 12119 129 12165
rect 175 12151 281 12165
rect 175 12119 287 12151
rect 333 12119 445 12165
rect 491 12119 620 12165
rect -58 12017 620 12119
rect -58 11965 281 12017
rect 333 11965 620 12017
rect -58 11944 620 11965
rect -58 11828 147 11944
rect -58 11782 -1 11828
rect 23 11782 147 11828
rect -58 11646 147 11782
rect -58 11600 -1 11646
rect 23 11600 147 11646
rect -58 11465 147 11600
rect -58 11419 -1 11465
rect 23 11419 147 11465
rect -58 11283 147 11419
rect -58 11237 -1 11283
rect 23 11237 147 11283
rect -58 11052 147 11237
rect 252 11828 367 11864
rect 252 11782 287 11828
rect 333 11782 367 11828
rect 252 11646 367 11782
rect 252 11633 287 11646
rect 333 11633 367 11646
rect 252 11477 285 11633
rect 337 11477 367 11633
rect 252 11465 367 11477
rect 252 11419 287 11465
rect 333 11419 367 11465
rect 252 11283 367 11419
rect 252 11237 287 11283
rect 333 11237 367 11283
rect 252 11200 367 11237
rect 472 11828 620 11944
rect 472 11782 513 11828
rect 559 11782 620 11828
rect 472 11646 620 11782
rect 472 11600 513 11646
rect 559 11600 620 11646
rect 472 11465 620 11600
rect 472 11419 513 11465
rect 559 11419 620 11465
rect 472 11283 620 11419
rect 472 11237 513 11283
rect 559 11237 620 11283
rect -58 11006 -1 11052
rect 23 11006 147 11052
rect -58 10871 147 11006
rect -58 10825 -1 10871
rect 23 10825 147 10871
rect -58 10690 147 10825
rect -58 10644 -1 10690
rect 23 10644 147 10690
rect -58 10508 147 10644
rect -58 10462 -1 10508
rect 23 10462 147 10508
rect -58 10425 147 10462
rect 252 11052 367 11089
rect 252 11006 287 11052
rect 333 11006 367 11052
rect 252 10871 367 11006
rect 252 10858 287 10871
rect 333 10858 367 10871
rect 252 10702 285 10858
rect 337 10702 367 10858
rect 252 10690 367 10702
rect 252 10644 287 10690
rect 333 10644 367 10690
rect 252 10508 367 10644
rect 252 10462 287 10508
rect 333 10462 367 10508
rect 252 10425 367 10462
rect 472 11052 620 11237
rect 472 11006 513 11052
rect 559 11006 620 11052
rect 472 10871 620 11006
rect 472 10825 513 10871
rect 559 10825 620 10871
rect 472 10690 620 10825
rect 472 10644 513 10690
rect 559 10644 620 10690
rect 472 10508 620 10644
rect 472 10462 513 10508
rect 559 10462 620 10508
rect 472 10425 620 10462
rect 159 10333 415 10344
rect 159 10287 170 10333
rect 404 10287 415 10333
rect 159 10276 415 10287
rect 58 9638 219 9650
rect 58 9482 70 9638
rect 122 9482 219 9638
rect 58 9470 219 9482
rect 397 9638 564 9650
rect 397 9482 500 9638
rect 552 9482 564 9638
rect 397 9470 564 9482
rect 70 8598 177 8610
rect 70 8442 82 8598
rect 134 8442 177 8598
rect 70 8045 177 8442
rect 114 7525 177 8045
rect 70 7248 177 7525
rect 433 7248 549 8610
rect 70 6919 141 7248
rect 219 7166 400 7178
rect 219 7010 290 7166
rect 342 7010 400 7166
rect 219 6995 400 7010
rect 479 6919 549 7248
rect 70 5557 184 6919
rect 443 5657 549 6919
rect 399 5567 549 5657
rect 399 5487 445 5567
rect 45 5465 445 5487
rect 45 5413 75 5465
rect 127 5413 445 5465
rect 45 5390 445 5413
rect -71 5306 71 5311
rect -71 5267 620 5306
rect -71 5260 368 5267
rect -71 5214 -23 5260
rect 23 5215 368 5260
rect 420 5215 620 5267
rect 23 5214 620 5215
rect -71 5172 620 5214
rect -71 5163 71 5172
rect 48 5059 565 5084
rect 48 5007 500 5059
rect 552 5007 565 5059
rect 48 4987 565 5007
rect 48 4915 141 4987
rect 48 3568 188 4915
rect 48 3553 192 3568
rect 443 3553 549 4907
rect 48 3060 141 3553
rect 219 3469 400 3483
rect 219 3459 287 3469
rect 333 3459 400 3469
rect 219 3407 286 3459
rect 338 3407 400 3459
rect 219 3348 400 3407
rect 219 3195 400 3268
rect 219 3143 284 3195
rect 336 3143 400 3195
rect 219 3132 400 3143
rect 272 3131 348 3132
rect 479 3060 549 3553
rect 48 1708 181 3060
rect 435 1710 549 3060
rect 364 1554 549 1710
rect -58 1415 620 1452
rect -58 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -58 1332 620 1369
rect -57 960 57 1332
rect 136 1227 404 1252
rect 136 1225 286 1227
rect 136 1179 230 1225
rect 276 1179 286 1225
rect 136 1175 286 1179
rect 338 1175 404 1227
rect 136 1155 404 1175
rect 549 1076 620 1332
rect -57 914 -23 960
rect 23 914 57 960
rect -57 797 57 914
rect 195 1064 303 1076
rect 195 908 226 1064
rect 278 908 303 1064
rect -57 271 57 500
rect 195 380 303 908
rect 446 960 620 1076
rect 446 914 480 960
rect 526 914 620 960
rect 446 797 620 914
rect 425 271 649 500
rect -58 147 649 271
rect -71 96 649 147
rect -71 50 -23 96
rect 23 50 135 96
rect 181 50 293 96
rect 339 50 451 96
rect 497 50 649 96
rect -71 -1 649 50
<< via1 >>
rect 281 12165 333 12203
rect 281 12151 287 12165
rect 287 12151 333 12165
rect 281 11965 333 12017
rect 285 11600 287 11633
rect 287 11600 333 11633
rect 333 11600 337 11633
rect 285 11477 337 11600
rect 285 10825 287 10858
rect 287 10825 333 10858
rect 333 10825 337 10858
rect 285 10702 337 10825
rect 70 9482 122 9638
rect 500 9482 552 9638
rect 82 8442 134 8598
rect 290 7164 342 7166
rect 290 7118 293 7164
rect 293 7118 339 7164
rect 339 7118 342 7164
rect 290 7010 342 7118
rect 75 5413 127 5465
rect 368 5215 420 5267
rect 500 5007 552 5059
rect 286 3423 287 3459
rect 287 3423 333 3459
rect 333 3423 338 3459
rect 286 3407 338 3423
rect 284 3192 336 3195
rect 284 3146 287 3192
rect 287 3146 333 3192
rect 333 3146 336 3192
rect 284 3143 336 3146
rect 286 1175 338 1227
rect 226 960 278 1064
rect 226 914 230 960
rect 230 914 276 960
rect 276 914 278 960
rect 226 908 278 914
<< metal2 >>
rect 68 11584 124 12225
rect 246 12205 374 12227
rect 246 12149 279 12205
rect 335 12149 374 12205
rect 246 12019 374 12149
rect 246 11963 279 12019
rect 335 11963 374 12019
rect 246 11944 374 11963
rect 273 11633 349 11645
rect 273 11584 285 11633
rect 68 11528 285 11584
rect 68 9650 124 11528
rect 273 11477 285 11528
rect 337 11477 349 11633
rect 273 11465 349 11477
rect 273 10858 349 10870
rect 273 10702 285 10858
rect 337 10808 349 10858
rect 498 10808 554 12225
rect 337 10752 554 10808
rect 337 10702 349 10752
rect 273 10690 349 10702
rect 498 9650 554 10752
rect 58 9638 134 9650
rect 58 9482 70 9638
rect 122 9482 134 9638
rect 58 9470 134 9482
rect 488 9638 564 9650
rect 488 9482 500 9638
rect 552 9482 564 9638
rect 488 9470 564 9482
rect 68 8610 124 9470
rect 68 8598 146 8610
rect 68 8442 82 8598
rect 134 8442 146 8598
rect 68 8430 146 8442
rect 278 7166 354 7178
rect 278 7010 290 7166
rect 342 7010 354 7166
rect 278 6998 354 7010
rect -28 5465 139 5477
rect -28 5413 75 5465
rect 127 5413 139 5465
rect -28 5401 139 5413
rect -28 -1 28 5401
rect 288 5397 344 6998
rect 221 5341 344 5397
rect 221 3655 277 5341
rect 356 5267 432 5279
rect 356 5256 368 5267
rect 420 5256 432 5267
rect 356 5096 366 5256
rect 422 5096 432 5256
rect 356 5086 432 5096
rect 498 5071 554 9470
rect 488 5059 564 5071
rect 488 5007 500 5059
rect 552 5007 564 5059
rect 488 4995 564 5007
rect 113 3599 277 3655
rect 113 3197 169 3599
rect 481 3483 573 4517
rect 250 3459 573 3483
rect 250 3407 286 3459
rect 338 3407 573 3459
rect 250 3386 573 3407
rect 272 3197 348 3207
rect 113 3195 348 3197
rect 113 3143 284 3195
rect 336 3143 348 3195
rect 113 3141 348 3143
rect 113 1076 169 3141
rect 272 3131 348 3141
rect 481 1853 573 3386
rect 274 1756 573 1853
rect 274 1227 350 1756
rect 274 1175 286 1227
rect 338 1175 350 1227
rect 274 1155 350 1175
rect 113 1064 290 1076
rect 113 908 226 1064
rect 278 908 290 1064
rect 113 896 290 908
rect 246 49 374 278
<< via2 >>
rect 279 12203 335 12205
rect 279 12151 281 12203
rect 281 12151 333 12203
rect 333 12151 335 12203
rect 279 12149 335 12151
rect 279 12017 335 12019
rect 279 11965 281 12017
rect 281 11965 333 12017
rect 333 11965 335 12017
rect 279 11963 335 11965
rect 366 5215 368 5256
rect 368 5215 420 5256
rect 420 5215 422 5256
rect 366 5096 422 5215
<< metal3 >>
rect -65 12205 929 12347
rect -65 12149 279 12205
rect 335 12149 929 12205
rect -65 12019 929 12149
rect -65 11963 279 12019
rect 335 11963 929 12019
rect -65 10538 929 11963
rect -1 5256 930 6638
rect -1 5096 366 5256
rect 422 5096 930 5256
rect -1 4657 930 5096
rect -1 4331 929 4546
rect -1 4009 929 4224
rect -1 3688 929 3903
rect -1 3366 929 3581
rect -1 2674 929 2889
rect -1 2352 929 2567
rect -1 2030 929 2245
rect -1 1708 929 1923
rect -1 1160 929 1602
rect -1 49 929 504
use M1_NWELL$$46277676_128x8m81  M1_NWELL$$46277676_128x8m81_0
timestamp 1666464484
transform 1 0 310 0 1 12142
box 0 0 1 1
use M1_NWELL$$47121452_128x8m81  M1_NWELL$$47121452_128x8m81_0
timestamp 1666464484
transform 1 0 237 0 1 1392
box 0 0 1 1
use M1_POLY24310590548731_128x8m81  M1_POLY24310590548731_128x8m81_0
timestamp 1666464484
transform 1 0 287 0 1 10310
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1666464484
transform 1 0 310 0 1 3446
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1666464484
transform 1 0 310 0 1 3169
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_2
timestamp 1666464484
transform 1 0 253 0 1 1202
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_3
timestamp 1666464484
transform 1 0 316 0 1 7141
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 5237
box 0 0 1 1
use M1_PSUB$$47122476_128x8m81  M1_PSUB$$47122476_128x8m81_0
timestamp 1666464484
transform 1 0 237 0 1 73
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1666464484
transform 1 0 311 0 1 10780
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_1
timestamp 1666464484
transform 1 0 311 0 1 11555
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_2
timestamp 1666464484
transform 1 0 96 0 1 9560
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_3
timestamp 1666464484
transform 1 0 108 0 1 8520
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_4
timestamp 1666464484
transform 1 0 252 0 1 986
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_5
timestamp 1666464484
transform 1 0 316 0 1 7088
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_6
timestamp 1666464484
transform 1 0 526 0 1 9560
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_0
timestamp 1666464484
transform 1 0 394 0 1 5241
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_1
timestamp 1666464484
transform 1 0 101 0 1 5439
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_2
timestamp 1666464484
transform 1 0 312 0 1 1201
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_3
timestamp 1666464484
transform 1 0 310 0 1 3169
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_4
timestamp 1666464484
transform 1 0 526 0 1 5033
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1666464484
transform 1 0 394 0 1 5176
box 0 0 1 1
use nmos_1p2$$47119404_128x8m81  nmos_1p2$$47119404_128x8m81_0
timestamp 1666464484
transform 1 0 281 0 -1 4915
box -119 -74 177 1434
use nmos_1p2$$47119404_128x8m81  nmos_1p2$$47119404_128x8m81_1
timestamp 1666464484
transform 1 0 281 0 -1 6919
box -119 -74 177 1434
use nmos_5p0431059054872_128x8m81  nmos_5p0431059054872_128x8m81_0
timestamp 1666464484
transform 1 0 52 0 1 383
box -88 -44 432 158
use pmos_1p2$$46889004_128x8m81  pmos_1p2$$46889004_128x8m81_0
timestamp 1666464484
transform 1 0 281 0 -1 3060
box -286 -142 343 1502
use pmos_5p0431059054871_128x8m81  pmos_5p0431059054871_128x8m81_0
timestamp 1666464484
transform 1 0 248 0 -1 10197
box -208 -120 328 1482
use pmos_5p0431059054871_128x8m81  pmos_5p0431059054871_128x8m81_1
timestamp 1666464484
transform 1 0 250 0 -1 8610
box -208 -120 328 1482
use via1_2_128x8m81  via1_2_128x8m81_0
timestamp 1666464484
transform 1 0 264 0 1 88
box -1 -1 93 128
use via1_R90_128x8m81  via1_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 378 1 0 3387
box 0 0 1 1
use via1_R90_128x8m81  via1_R90_128x8m81_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
use via1_R90_128x8m81  via1_R90_128x8m81_2
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_128x8m81  via2_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_128x8m81  via2_R90_128x8m81_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
<< labels >>
rlabel metal3 s 279 91 279 91 4 vss
port 1 nsew
rlabel metal3 s 318 12094 318 12094 4 vdd
port 2 nsew
rlabel metal3 s 303 5255 303 5255 4 vss
port 1 nsew
rlabel metal2 s 518 11931 518 11931 4 b
port 3 nsew
rlabel metal2 s 105 11931 105 11931 4 bb
port 4 nsew
rlabel metal2 s 0 304 0 304 4 db
port 5 nsew
rlabel metal2 s 285 1222 285 1222 4 ypass
port 6 nsew
rlabel metal1 s 492 1805 492 1805 4 d
port 7 nsew
rlabel metal1 s 259 10292 259 10292 4 pcb
port 8 nsew
rlabel metal1 s 318 1356 318 1356 4 vdd
port 2 nsew
<< properties >>
string GDS_END 302300
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 293038
string path 0.000 27.385 0.000 -0.005 
<< end >>
