magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 2360 686
<< polysilicon >>
rect -31 544 89 618
rect 193 544 313 618
rect 417 544 537 618
rect 641 544 761 618
rect 865 544 985 618
rect 1089 544 1209 618
rect 1313 544 1433 618
rect 1537 544 1657 618
rect 1761 544 1881 618
rect 1985 544 2105 618
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 641 -74 761 -1
rect 865 -74 985 -1
rect 1089 -74 1209 -1
rect 1313 -74 1433 -1
rect 1537 -74 1657 -1
rect 1761 -74 1881 -1
rect 1985 -74 2105 -1
use pmos_5p04310590878128_256x8m81  pmos_5p04310590878128_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 2344 664
<< properties >>
string GDS_END 349012
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 347546
<< end >>
