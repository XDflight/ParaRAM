magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 4118 1094
<< pwell >>
rect -86 -86 4118 453
<< mvnmos >>
rect 124 146 244 304
rect 348 146 468 304
rect 720 215 840 333
rect 944 215 1064 333
rect 1168 215 1288 333
rect 1336 215 1456 333
rect 1568 215 1688 333
rect 1736 215 1856 333
rect 1960 215 2080 333
rect 2220 183 2340 333
rect 2816 183 2936 333
rect 3076 215 3196 333
rect 3336 183 3456 333
rect 3704 69 3824 333
<< mvpmos >>
rect 124 573 224 849
rect 328 573 428 849
rect 720 573 820 773
rect 924 573 1024 773
rect 1128 573 1228 773
rect 1276 573 1376 773
rect 1568 573 1668 773
rect 1816 651 1916 851
rect 2248 573 2348 773
rect 2488 573 2588 793
rect 2836 633 2936 853
rect 3096 579 3196 779
rect 3344 579 3444 799
rect 3704 573 3804 939
<< mvndiff >>
rect 36 291 124 304
rect 36 245 49 291
rect 95 245 124 291
rect 36 146 124 245
rect 244 205 348 304
rect 244 159 273 205
rect 319 159 348 205
rect 244 146 348 159
rect 468 291 556 304
rect 468 245 497 291
rect 543 245 556 291
rect 468 146 556 245
rect 632 274 720 333
rect 632 228 645 274
rect 691 228 720 274
rect 632 215 720 228
rect 840 320 944 333
rect 840 274 869 320
rect 915 274 944 320
rect 840 215 944 274
rect 1064 320 1168 333
rect 1064 274 1093 320
rect 1139 274 1168 320
rect 1064 215 1168 274
rect 1288 215 1336 333
rect 1456 274 1568 333
rect 1456 228 1485 274
rect 1531 228 1568 274
rect 1456 215 1568 228
rect 1688 215 1736 333
rect 1856 320 1960 333
rect 1856 274 1885 320
rect 1931 274 1960 320
rect 1856 215 1960 274
rect 2080 320 2220 333
rect 2080 274 2145 320
rect 2191 274 2220 320
rect 2080 215 2220 274
rect 2140 183 2220 215
rect 2340 298 2428 333
rect 2340 252 2369 298
rect 2415 252 2428 298
rect 2340 183 2428 252
rect 2725 320 2816 333
rect 2725 274 2738 320
rect 2784 274 2816 320
rect 2725 183 2816 274
rect 2936 215 3076 333
rect 3196 273 3336 333
rect 3196 227 3261 273
rect 3307 227 3336 273
rect 3196 215 3336 227
rect 2936 183 3016 215
rect 3256 183 3336 215
rect 3456 320 3544 333
rect 3456 274 3485 320
rect 3531 274 3544 320
rect 3456 183 3544 274
rect 3616 320 3704 333
rect 3616 180 3629 320
rect 3675 180 3704 320
rect 3616 69 3704 180
rect 3824 222 3912 333
rect 3824 82 3853 222
rect 3899 82 3912 222
rect 3824 69 3912 82
<< mvpdiff >>
rect 36 726 124 849
rect 36 586 49 726
rect 95 586 124 726
rect 36 573 124 586
rect 224 836 328 849
rect 224 696 253 836
rect 299 696 328 836
rect 224 573 328 696
rect 428 726 516 849
rect 428 586 457 726
rect 503 586 516 726
rect 428 573 516 586
rect 588 838 660 851
rect 588 792 601 838
rect 647 792 660 838
rect 588 773 660 792
rect 1436 932 1508 945
rect 1436 792 1449 932
rect 1495 792 1508 932
rect 1436 773 1508 792
rect 1736 773 1816 851
rect 588 573 720 773
rect 820 643 924 773
rect 820 597 849 643
rect 895 597 924 643
rect 820 573 924 597
rect 1024 632 1128 773
rect 1024 586 1053 632
rect 1099 586 1128 632
rect 1024 573 1128 586
rect 1228 573 1276 773
rect 1376 573 1568 773
rect 1668 651 1816 773
rect 1916 838 2004 851
rect 1916 792 1945 838
rect 1991 792 2004 838
rect 1916 651 2004 792
rect 2748 840 2836 853
rect 2748 794 2761 840
rect 2807 794 2836 840
rect 2408 773 2488 793
rect 1668 632 1756 651
rect 1668 586 1697 632
rect 1743 586 1756 632
rect 1668 573 1756 586
rect 2160 632 2248 773
rect 2160 586 2173 632
rect 2219 586 2248 632
rect 2160 573 2248 586
rect 2348 726 2488 773
rect 2348 586 2377 726
rect 2423 586 2488 726
rect 2348 573 2488 586
rect 2588 632 2676 793
rect 2748 633 2836 794
rect 2936 779 3016 853
rect 3256 786 3344 799
rect 3256 779 3269 786
rect 2936 638 3096 779
rect 2936 633 3021 638
rect 2588 586 2617 632
rect 2663 586 2676 632
rect 2588 573 2676 586
rect 3008 592 3021 633
rect 3067 592 3096 638
rect 3008 579 3096 592
rect 3196 646 3269 779
rect 3315 646 3344 786
rect 3196 579 3344 646
rect 3444 732 3532 799
rect 3444 592 3473 732
rect 3519 592 3532 732
rect 3444 579 3532 592
rect 3616 726 3704 939
rect 3616 586 3629 726
rect 3675 586 3704 726
rect 3616 573 3704 586
rect 3804 926 3892 939
rect 3804 786 3833 926
rect 3879 786 3892 926
rect 3804 573 3892 786
<< mvndiffc >>
rect 49 245 95 291
rect 273 159 319 205
rect 497 245 543 291
rect 645 228 691 274
rect 869 274 915 320
rect 1093 274 1139 320
rect 1485 228 1531 274
rect 1885 274 1931 320
rect 2145 274 2191 320
rect 2369 252 2415 298
rect 2738 274 2784 320
rect 3261 227 3307 273
rect 3485 274 3531 320
rect 3629 180 3675 320
rect 3853 82 3899 222
<< mvpdiffc >>
rect 49 586 95 726
rect 253 696 299 836
rect 457 586 503 726
rect 601 792 647 838
rect 1449 792 1495 932
rect 849 597 895 643
rect 1053 586 1099 632
rect 1945 792 1991 838
rect 2761 794 2807 840
rect 1697 586 1743 632
rect 2173 586 2219 632
rect 2377 586 2423 726
rect 2617 586 2663 632
rect 3021 592 3067 638
rect 3269 646 3315 786
rect 3473 592 3519 732
rect 3629 586 3675 726
rect 3833 786 3879 926
<< polysilicon >>
rect 328 911 1024 951
rect 124 849 224 893
rect 328 849 428 911
rect 720 773 820 817
rect 924 773 1024 911
rect 1128 852 1228 865
rect 1128 806 1141 852
rect 1187 806 1228 852
rect 1128 773 1228 806
rect 1276 773 1376 817
rect 1816 913 2936 953
rect 3704 939 3804 983
rect 1816 851 1916 913
rect 2248 852 2348 865
rect 2836 853 2936 913
rect 1568 773 1668 817
rect 2248 806 2261 852
rect 2307 806 2348 852
rect 2248 773 2348 806
rect 2488 793 2588 837
rect 1816 607 1916 651
rect 124 400 224 573
rect 124 354 137 400
rect 183 354 224 400
rect 328 383 428 573
rect 328 364 361 383
rect 124 348 224 354
rect 124 304 244 348
rect 348 337 361 364
rect 407 364 428 383
rect 720 523 820 573
rect 924 529 1024 573
rect 720 477 733 523
rect 779 477 820 523
rect 1128 481 1228 573
rect 720 377 820 477
rect 944 441 1228 481
rect 1276 540 1376 573
rect 1276 494 1317 540
rect 1363 494 1376 540
rect 407 337 468 364
rect 348 304 468 337
rect 720 333 840 377
rect 944 333 1064 441
rect 1276 425 1376 494
rect 1168 333 1288 377
rect 1336 333 1456 425
rect 1568 412 1668 573
rect 1568 366 1581 412
rect 1627 377 1668 412
rect 1816 377 1856 607
rect 3096 779 3196 823
rect 3344 799 3444 843
rect 2248 529 2348 573
rect 2248 377 2340 529
rect 1627 366 1688 377
rect 1568 333 1688 366
rect 1736 333 1856 377
rect 1960 333 2080 377
rect 2220 333 2340 377
rect 720 171 840 215
rect 944 171 1064 215
rect 124 102 244 146
rect 348 86 468 146
rect 1168 86 1288 215
rect 1336 171 1456 215
rect 1568 171 1688 215
rect 1736 171 1856 215
rect 1960 86 2080 215
rect 2220 139 2340 183
rect 2488 86 2588 573
rect 2836 510 2936 633
rect 2836 464 2849 510
rect 2895 464 2936 510
rect 2836 377 2936 464
rect 3096 443 3196 579
rect 3096 397 3137 443
rect 3183 397 3196 443
rect 3096 377 3196 397
rect 3344 546 3444 579
rect 3344 500 3357 546
rect 3403 500 3444 546
rect 3344 377 3444 500
rect 3704 465 3804 573
rect 3524 452 3804 465
rect 3524 406 3537 452
rect 3583 406 3804 452
rect 3524 393 3804 406
rect 3704 377 3804 393
rect 2816 333 2936 377
rect 3076 333 3196 377
rect 3336 333 3456 377
rect 3704 333 3824 377
rect 2816 139 2936 183
rect 3076 171 3196 215
rect 3336 139 3456 183
rect 348 46 2588 86
rect 3704 25 3824 69
<< polycontact >>
rect 1141 806 1187 852
rect 2261 806 2307 852
rect 137 354 183 400
rect 361 337 407 383
rect 733 477 779 523
rect 1317 494 1363 540
rect 1581 366 1627 412
rect 2849 464 2895 510
rect 3137 397 3183 443
rect 3357 500 3403 546
rect 3537 406 3583 452
<< metal1 >>
rect 0 932 4032 1098
rect 0 918 1449 932
rect 253 836 299 918
rect 49 726 95 737
rect 601 838 647 918
rect 601 781 647 792
rect 1130 806 1141 852
rect 1187 806 1198 852
rect 253 685 299 696
rect 457 735 503 737
rect 1130 735 1198 806
rect 1495 926 4032 932
rect 1495 918 3833 926
rect 1449 781 1495 792
rect 1945 838 1991 918
rect 1945 781 1991 792
rect 2261 852 2307 863
rect 2261 735 2307 806
rect 2761 840 2807 918
rect 2761 783 2807 794
rect 3269 786 3315 918
rect 2826 737 3223 741
rect 457 726 2307 735
rect 95 586 407 621
rect 49 575 407 586
rect 126 400 306 430
rect 126 354 137 400
rect 183 354 306 400
rect 361 383 407 575
rect 361 308 407 337
rect 49 291 407 308
rect 95 262 407 291
rect 503 689 2307 726
rect 2377 726 3223 737
rect 503 586 543 689
rect 457 291 543 586
rect 610 597 849 643
rect 895 597 906 643
rect 1053 632 1099 643
rect 610 420 656 597
rect 702 523 910 542
rect 702 477 733 523
rect 779 477 910 523
rect 702 466 910 477
rect 610 374 783 420
rect 49 234 95 245
rect 457 245 497 291
rect 737 331 783 374
rect 1053 412 1099 586
rect 1697 632 1743 643
rect 1697 540 1743 586
rect 2173 632 2219 643
rect 2173 540 2219 586
rect 1306 494 1317 540
rect 1363 494 2219 540
rect 2423 695 3223 726
rect 2423 691 2845 695
rect 3021 643 3067 649
rect 1053 366 1581 412
rect 1627 366 1638 412
rect 737 320 915 331
rect 457 234 543 245
rect 645 274 691 285
rect 737 274 869 320
rect 737 263 915 274
rect 1053 320 1139 366
rect 1053 274 1093 320
rect 1885 320 1931 494
rect 2377 401 2423 586
rect 2617 638 3067 643
rect 2617 632 3021 638
rect 2663 597 3021 632
rect 2663 586 2784 597
rect 2617 575 2784 586
rect 3021 581 3067 592
rect 1053 263 1139 274
rect 1485 274 1531 285
rect 273 205 319 216
rect 273 90 319 159
rect 645 90 691 228
rect 1885 263 1931 274
rect 2145 355 2423 401
rect 2145 320 2191 355
rect 2738 320 2784 575
rect 3177 546 3223 695
rect 3879 918 4032 926
rect 3833 775 3879 786
rect 3269 635 3315 646
rect 3473 732 3519 743
rect 2830 510 2995 542
rect 2830 464 2849 510
rect 2895 464 2995 510
rect 3177 500 3357 546
rect 3403 500 3414 546
rect 2830 453 2995 464
rect 3473 463 3519 592
rect 3629 726 3675 737
rect 3473 454 3583 463
rect 3137 452 3583 454
rect 3137 443 3537 452
rect 3183 406 3537 443
rect 3183 397 3583 406
rect 3137 395 3583 397
rect 3137 386 3531 395
rect 2145 263 2191 274
rect 2369 298 2738 309
rect 2415 274 2738 298
rect 3485 320 3531 386
rect 2415 252 2784 274
rect 2369 241 2784 252
rect 3261 273 3307 284
rect 1485 90 1531 228
rect 3629 320 3675 586
rect 3485 263 3531 274
rect 3261 90 3307 227
rect 3614 180 3629 318
rect 3614 169 3675 180
rect 3853 222 3899 233
rect 0 82 3853 90
rect 3899 82 4032 90
rect 0 -90 4032 82
<< labels >>
flabel metal1 s 126 354 306 430 0 FreeSans 200 0 0 0 CLKN
port 3 nsew clock input
flabel metal1 s 702 466 910 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3629 318 3675 737 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 2830 453 2995 542 0 FreeSans 200 0 0 0 SETN
port 2 nsew default input
flabel metal1 s 0 918 4032 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1485 284 1531 285 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3614 169 3675 318 1 Q
port 4 nsew default output
rlabel metal1 s 3833 783 3879 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3269 783 3315 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2761 783 2807 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1945 783 1991 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1449 783 1495 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 601 783 647 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 253 783 299 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3833 781 3879 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3269 781 3315 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1945 781 1991 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1449 781 1495 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 601 781 647 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 253 781 299 783 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3833 775 3879 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3269 775 3315 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 253 775 299 781 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3269 685 3315 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 253 685 299 775 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3269 635 3315 685 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 645 284 691 285 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3261 233 3307 284 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1485 233 1531 284 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 645 233 691 284 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3853 216 3899 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3261 216 3307 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1485 216 1531 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 645 216 691 233 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3853 90 3899 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3261 90 3307 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1485 90 1531 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 645 90 691 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4032 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 1008
string GDS_END 550180
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 541678
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
