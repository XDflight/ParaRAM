magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -236 510 236 515
rect -236 482 -231 510
rect -203 482 -169 510
rect -141 482 -107 510
rect -79 482 -45 510
rect -17 482 17 510
rect 45 482 79 510
rect 107 482 141 510
rect 169 482 203 510
rect 231 482 236 510
rect -236 448 236 482
rect -236 420 -231 448
rect -203 420 -169 448
rect -141 420 -107 448
rect -79 420 -45 448
rect -17 420 17 448
rect 45 420 79 448
rect 107 420 141 448
rect 169 420 203 448
rect 231 420 236 448
rect -236 386 236 420
rect -236 358 -231 386
rect -203 358 -169 386
rect -141 358 -107 386
rect -79 358 -45 386
rect -17 358 17 386
rect 45 358 79 386
rect 107 358 141 386
rect 169 358 203 386
rect 231 358 236 386
rect -236 324 236 358
rect -236 296 -231 324
rect -203 296 -169 324
rect -141 296 -107 324
rect -79 296 -45 324
rect -17 296 17 324
rect 45 296 79 324
rect 107 296 141 324
rect 169 296 203 324
rect 231 296 236 324
rect -236 262 236 296
rect -236 234 -231 262
rect -203 234 -169 262
rect -141 234 -107 262
rect -79 234 -45 262
rect -17 234 17 262
rect 45 234 79 262
rect 107 234 141 262
rect 169 234 203 262
rect 231 234 236 262
rect -236 200 236 234
rect -236 172 -231 200
rect -203 172 -169 200
rect -141 172 -107 200
rect -79 172 -45 200
rect -17 172 17 200
rect 45 172 79 200
rect 107 172 141 200
rect 169 172 203 200
rect 231 172 236 200
rect -236 138 236 172
rect -236 110 -231 138
rect -203 110 -169 138
rect -141 110 -107 138
rect -79 110 -45 138
rect -17 110 17 138
rect 45 110 79 138
rect 107 110 141 138
rect 169 110 203 138
rect 231 110 236 138
rect -236 76 236 110
rect -236 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 236 76
rect -236 14 236 48
rect -236 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 236 14
rect -236 -48 236 -14
rect -236 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 236 -48
rect -236 -110 236 -76
rect -236 -138 -231 -110
rect -203 -138 -169 -110
rect -141 -138 -107 -110
rect -79 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 79 -110
rect 107 -138 141 -110
rect 169 -138 203 -110
rect 231 -138 236 -110
rect -236 -172 236 -138
rect -236 -200 -231 -172
rect -203 -200 -169 -172
rect -141 -200 -107 -172
rect -79 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 79 -172
rect 107 -200 141 -172
rect 169 -200 203 -172
rect 231 -200 236 -172
rect -236 -234 236 -200
rect -236 -262 -231 -234
rect -203 -262 -169 -234
rect -141 -262 -107 -234
rect -79 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 79 -234
rect 107 -262 141 -234
rect 169 -262 203 -234
rect 231 -262 236 -234
rect -236 -296 236 -262
rect -236 -324 -231 -296
rect -203 -324 -169 -296
rect -141 -324 -107 -296
rect -79 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 79 -296
rect 107 -324 141 -296
rect 169 -324 203 -296
rect 231 -324 236 -296
rect -236 -358 236 -324
rect -236 -386 -231 -358
rect -203 -386 -169 -358
rect -141 -386 -107 -358
rect -79 -386 -45 -358
rect -17 -386 17 -358
rect 45 -386 79 -358
rect 107 -386 141 -358
rect 169 -386 203 -358
rect 231 -386 236 -358
rect -236 -420 236 -386
rect -236 -448 -231 -420
rect -203 -448 -169 -420
rect -141 -448 -107 -420
rect -79 -448 -45 -420
rect -17 -448 17 -420
rect 45 -448 79 -420
rect 107 -448 141 -420
rect 169 -448 203 -420
rect 231 -448 236 -420
rect -236 -482 236 -448
rect -236 -510 -231 -482
rect -203 -510 -169 -482
rect -141 -510 -107 -482
rect -79 -510 -45 -482
rect -17 -510 17 -482
rect 45 -510 79 -482
rect 107 -510 141 -482
rect 169 -510 203 -482
rect 231 -510 236 -482
rect -236 -515 236 -510
<< via2 >>
rect -231 482 -203 510
rect -169 482 -141 510
rect -107 482 -79 510
rect -45 482 -17 510
rect 17 482 45 510
rect 79 482 107 510
rect 141 482 169 510
rect 203 482 231 510
rect -231 420 -203 448
rect -169 420 -141 448
rect -107 420 -79 448
rect -45 420 -17 448
rect 17 420 45 448
rect 79 420 107 448
rect 141 420 169 448
rect 203 420 231 448
rect -231 358 -203 386
rect -169 358 -141 386
rect -107 358 -79 386
rect -45 358 -17 386
rect 17 358 45 386
rect 79 358 107 386
rect 141 358 169 386
rect 203 358 231 386
rect -231 296 -203 324
rect -169 296 -141 324
rect -107 296 -79 324
rect -45 296 -17 324
rect 17 296 45 324
rect 79 296 107 324
rect 141 296 169 324
rect 203 296 231 324
rect -231 234 -203 262
rect -169 234 -141 262
rect -107 234 -79 262
rect -45 234 -17 262
rect 17 234 45 262
rect 79 234 107 262
rect 141 234 169 262
rect 203 234 231 262
rect -231 172 -203 200
rect -169 172 -141 200
rect -107 172 -79 200
rect -45 172 -17 200
rect 17 172 45 200
rect 79 172 107 200
rect 141 172 169 200
rect 203 172 231 200
rect -231 110 -203 138
rect -169 110 -141 138
rect -107 110 -79 138
rect -45 110 -17 138
rect 17 110 45 138
rect 79 110 107 138
rect 141 110 169 138
rect 203 110 231 138
rect -231 48 -203 76
rect -169 48 -141 76
rect -107 48 -79 76
rect -45 48 -17 76
rect 17 48 45 76
rect 79 48 107 76
rect 141 48 169 76
rect 203 48 231 76
rect -231 -14 -203 14
rect -169 -14 -141 14
rect -107 -14 -79 14
rect -45 -14 -17 14
rect 17 -14 45 14
rect 79 -14 107 14
rect 141 -14 169 14
rect 203 -14 231 14
rect -231 -76 -203 -48
rect -169 -76 -141 -48
rect -107 -76 -79 -48
rect -45 -76 -17 -48
rect 17 -76 45 -48
rect 79 -76 107 -48
rect 141 -76 169 -48
rect 203 -76 231 -48
rect -231 -138 -203 -110
rect -169 -138 -141 -110
rect -107 -138 -79 -110
rect -45 -138 -17 -110
rect 17 -138 45 -110
rect 79 -138 107 -110
rect 141 -138 169 -110
rect 203 -138 231 -110
rect -231 -200 -203 -172
rect -169 -200 -141 -172
rect -107 -200 -79 -172
rect -45 -200 -17 -172
rect 17 -200 45 -172
rect 79 -200 107 -172
rect 141 -200 169 -172
rect 203 -200 231 -172
rect -231 -262 -203 -234
rect -169 -262 -141 -234
rect -107 -262 -79 -234
rect -45 -262 -17 -234
rect 17 -262 45 -234
rect 79 -262 107 -234
rect 141 -262 169 -234
rect 203 -262 231 -234
rect -231 -324 -203 -296
rect -169 -324 -141 -296
rect -107 -324 -79 -296
rect -45 -324 -17 -296
rect 17 -324 45 -296
rect 79 -324 107 -296
rect 141 -324 169 -296
rect 203 -324 231 -296
rect -231 -386 -203 -358
rect -169 -386 -141 -358
rect -107 -386 -79 -358
rect -45 -386 -17 -358
rect 17 -386 45 -358
rect 79 -386 107 -358
rect 141 -386 169 -358
rect 203 -386 231 -358
rect -231 -448 -203 -420
rect -169 -448 -141 -420
rect -107 -448 -79 -420
rect -45 -448 -17 -420
rect 17 -448 45 -420
rect 79 -448 107 -420
rect 141 -448 169 -420
rect 203 -448 231 -420
rect -231 -510 -203 -482
rect -169 -510 -141 -482
rect -107 -510 -79 -482
rect -45 -510 -17 -482
rect 17 -510 45 -482
rect 79 -510 107 -482
rect 141 -510 169 -482
rect 203 -510 231 -482
<< metal3 >>
rect -236 510 236 515
rect -236 482 -231 510
rect -203 482 -169 510
rect -141 482 -107 510
rect -79 482 -45 510
rect -17 482 17 510
rect 45 482 79 510
rect 107 482 141 510
rect 169 482 203 510
rect 231 482 236 510
rect -236 448 236 482
rect -236 420 -231 448
rect -203 420 -169 448
rect -141 420 -107 448
rect -79 420 -45 448
rect -17 420 17 448
rect 45 420 79 448
rect 107 420 141 448
rect 169 420 203 448
rect 231 420 236 448
rect -236 386 236 420
rect -236 358 -231 386
rect -203 358 -169 386
rect -141 358 -107 386
rect -79 358 -45 386
rect -17 358 17 386
rect 45 358 79 386
rect 107 358 141 386
rect 169 358 203 386
rect 231 358 236 386
rect -236 324 236 358
rect -236 296 -231 324
rect -203 296 -169 324
rect -141 296 -107 324
rect -79 296 -45 324
rect -17 296 17 324
rect 45 296 79 324
rect 107 296 141 324
rect 169 296 203 324
rect 231 296 236 324
rect -236 262 236 296
rect -236 234 -231 262
rect -203 234 -169 262
rect -141 234 -107 262
rect -79 234 -45 262
rect -17 234 17 262
rect 45 234 79 262
rect 107 234 141 262
rect 169 234 203 262
rect 231 234 236 262
rect -236 200 236 234
rect -236 172 -231 200
rect -203 172 -169 200
rect -141 172 -107 200
rect -79 172 -45 200
rect -17 172 17 200
rect 45 172 79 200
rect 107 172 141 200
rect 169 172 203 200
rect 231 172 236 200
rect -236 138 236 172
rect -236 110 -231 138
rect -203 110 -169 138
rect -141 110 -107 138
rect -79 110 -45 138
rect -17 110 17 138
rect 45 110 79 138
rect 107 110 141 138
rect 169 110 203 138
rect 231 110 236 138
rect -236 76 236 110
rect -236 48 -231 76
rect -203 48 -169 76
rect -141 48 -107 76
rect -79 48 -45 76
rect -17 48 17 76
rect 45 48 79 76
rect 107 48 141 76
rect 169 48 203 76
rect 231 48 236 76
rect -236 14 236 48
rect -236 -14 -231 14
rect -203 -14 -169 14
rect -141 -14 -107 14
rect -79 -14 -45 14
rect -17 -14 17 14
rect 45 -14 79 14
rect 107 -14 141 14
rect 169 -14 203 14
rect 231 -14 236 14
rect -236 -48 236 -14
rect -236 -76 -231 -48
rect -203 -76 -169 -48
rect -141 -76 -107 -48
rect -79 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 79 -48
rect 107 -76 141 -48
rect 169 -76 203 -48
rect 231 -76 236 -48
rect -236 -110 236 -76
rect -236 -138 -231 -110
rect -203 -138 -169 -110
rect -141 -138 -107 -110
rect -79 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 79 -110
rect 107 -138 141 -110
rect 169 -138 203 -110
rect 231 -138 236 -110
rect -236 -172 236 -138
rect -236 -200 -231 -172
rect -203 -200 -169 -172
rect -141 -200 -107 -172
rect -79 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 79 -172
rect 107 -200 141 -172
rect 169 -200 203 -172
rect 231 -200 236 -172
rect -236 -234 236 -200
rect -236 -262 -231 -234
rect -203 -262 -169 -234
rect -141 -262 -107 -234
rect -79 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 79 -234
rect 107 -262 141 -234
rect 169 -262 203 -234
rect 231 -262 236 -234
rect -236 -296 236 -262
rect -236 -324 -231 -296
rect -203 -324 -169 -296
rect -141 -324 -107 -296
rect -79 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 79 -296
rect 107 -324 141 -296
rect 169 -324 203 -296
rect 231 -324 236 -296
rect -236 -358 236 -324
rect -236 -386 -231 -358
rect -203 -386 -169 -358
rect -141 -386 -107 -358
rect -79 -386 -45 -358
rect -17 -386 17 -358
rect 45 -386 79 -358
rect 107 -386 141 -358
rect 169 -386 203 -358
rect 231 -386 236 -358
rect -236 -420 236 -386
rect -236 -448 -231 -420
rect -203 -448 -169 -420
rect -141 -448 -107 -420
rect -79 -448 -45 -420
rect -17 -448 17 -420
rect 45 -448 79 -420
rect 107 -448 141 -420
rect 169 -448 203 -420
rect 231 -448 236 -420
rect -236 -482 236 -448
rect -236 -510 -231 -482
rect -203 -510 -169 -482
rect -141 -510 -107 -482
rect -79 -510 -45 -482
rect -17 -510 17 -482
rect 45 -510 79 -482
rect 107 -510 141 -482
rect 169 -510 203 -482
rect 231 -510 236 -482
rect -236 -515 236 -510
<< properties >>
string GDS_END 734978
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 726142
<< end >>
