magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 2886 870
<< pwell >>
rect -86 -86 2886 352
<< mvnmos >>
rect 131 68 251 228
rect 299 68 419 228
rect 577 68 697 228
rect 759 68 879 228
rect 1071 68 1191 228
rect 1275 68 1395 228
rect 1499 68 1619 228
rect 1683 68 1803 228
rect 1910 68 2030 228
rect 2094 68 2214 228
rect 2318 68 2438 228
rect 2502 68 2622 228
<< mvpmos >>
rect 131 472 231 716
rect 335 472 435 716
rect 539 472 639 716
rect 743 472 843 716
rect 1091 472 1191 716
rect 1295 472 1395 716
rect 1499 472 1599 716
rect 1703 472 1803 716
rect 1910 472 2010 716
rect 2114 472 2214 716
rect 2318 472 2418 716
rect 2522 472 2622 716
<< mvndiff >>
rect 43 194 131 228
rect 43 148 56 194
rect 102 148 131 194
rect 43 68 131 148
rect 251 68 299 228
rect 419 127 577 228
rect 419 81 502 127
rect 548 81 577 127
rect 419 68 577 81
rect 697 68 759 228
rect 879 215 1071 228
rect 879 169 996 215
rect 1042 169 1071 215
rect 879 68 1071 169
rect 1191 68 1275 228
rect 1395 127 1499 228
rect 1395 81 1424 127
rect 1470 81 1499 127
rect 1395 68 1499 81
rect 1619 68 1683 228
rect 1803 215 1910 228
rect 1803 169 1832 215
rect 1878 169 1910 215
rect 1803 68 1910 169
rect 2030 68 2094 228
rect 2214 127 2318 228
rect 2214 81 2243 127
rect 2289 81 2318 127
rect 2214 68 2318 81
rect 2438 68 2502 228
rect 2622 171 2710 228
rect 2622 125 2651 171
rect 2697 125 2710 171
rect 2622 68 2710 125
<< mvpdiff >>
rect 43 665 131 716
rect 43 525 56 665
rect 102 525 131 665
rect 43 472 131 525
rect 231 665 335 716
rect 231 525 260 665
rect 306 525 335 665
rect 231 472 335 525
rect 435 665 539 716
rect 435 619 464 665
rect 510 619 539 665
rect 435 472 539 619
rect 639 665 743 716
rect 639 525 668 665
rect 714 525 743 665
rect 639 472 743 525
rect 843 665 931 716
rect 843 619 872 665
rect 918 619 931 665
rect 843 472 931 619
rect 1003 678 1091 716
rect 1003 632 1016 678
rect 1062 632 1091 678
rect 1003 472 1091 632
rect 1191 552 1295 716
rect 1191 506 1220 552
rect 1266 506 1295 552
rect 1191 472 1295 506
rect 1395 678 1499 716
rect 1395 632 1424 678
rect 1470 632 1499 678
rect 1395 472 1499 632
rect 1599 552 1703 716
rect 1599 506 1628 552
rect 1674 506 1703 552
rect 1599 472 1703 506
rect 1803 678 1910 716
rect 1803 632 1832 678
rect 1878 632 1910 678
rect 1803 472 1910 632
rect 2010 534 2114 716
rect 2010 488 2039 534
rect 2085 488 2114 534
rect 2010 472 2114 488
rect 2214 678 2318 716
rect 2214 632 2243 678
rect 2289 632 2318 678
rect 2214 472 2318 632
rect 2418 534 2522 716
rect 2418 488 2447 534
rect 2493 488 2522 534
rect 2418 472 2522 488
rect 2622 678 2710 716
rect 2622 632 2651 678
rect 2697 632 2710 678
rect 2622 472 2710 632
<< mvndiffc >>
rect 56 148 102 194
rect 502 81 548 127
rect 996 169 1042 215
rect 1424 81 1470 127
rect 1832 169 1878 215
rect 2243 81 2289 127
rect 2651 125 2697 171
<< mvpdiffc >>
rect 56 525 102 665
rect 260 525 306 665
rect 464 619 510 665
rect 668 525 714 665
rect 872 619 918 665
rect 1016 632 1062 678
rect 1220 506 1266 552
rect 1424 632 1470 678
rect 1628 506 1674 552
rect 1832 632 1878 678
rect 2039 488 2085 534
rect 2243 632 2289 678
rect 2447 488 2493 534
rect 2651 632 2697 678
<< polysilicon >>
rect 131 716 231 760
rect 335 716 435 760
rect 539 716 639 760
rect 743 716 843 760
rect 1091 716 1191 760
rect 1295 716 1395 760
rect 1499 716 1599 760
rect 1703 716 1803 760
rect 1910 716 2010 760
rect 2114 716 2214 760
rect 2318 716 2418 760
rect 2522 716 2622 760
rect 131 439 231 472
rect 131 393 155 439
rect 201 393 231 439
rect 131 288 231 393
rect 335 332 435 472
rect 539 351 639 472
rect 743 439 843 472
rect 743 393 764 439
rect 810 393 843 439
rect 743 380 843 393
rect 539 332 697 351
rect 335 324 697 332
rect 299 314 697 324
rect 299 307 614 314
rect 131 228 251 288
rect 299 261 312 307
rect 358 292 614 307
rect 358 261 419 292
rect 299 228 419 261
rect 577 268 614 292
rect 660 268 697 314
rect 577 228 697 268
rect 759 276 843 380
rect 1091 311 1191 472
rect 1295 439 1395 472
rect 1295 393 1308 439
rect 1354 393 1395 439
rect 1295 333 1395 393
rect 1499 333 1599 472
rect 1703 406 1803 472
rect 1295 332 1599 333
rect 1091 288 1132 311
rect 759 228 879 276
rect 1071 265 1132 288
rect 1178 265 1191 311
rect 1071 228 1191 265
rect 1275 293 1599 332
rect 1275 228 1395 293
rect 1499 288 1599 293
rect 1683 393 1803 406
rect 1683 347 1696 393
rect 1742 347 1803 393
rect 1499 228 1619 288
rect 1683 228 1803 347
rect 1910 439 2010 472
rect 1910 393 1951 439
rect 1997 393 2010 439
rect 1910 288 2010 393
rect 2114 332 2214 472
rect 2318 332 2418 472
rect 2114 313 2418 332
rect 2114 288 2144 313
rect 1910 228 2030 288
rect 2094 267 2144 288
rect 2190 292 2344 313
rect 2190 267 2214 292
rect 2094 228 2214 267
rect 2318 267 2344 292
rect 2390 288 2418 313
rect 2522 403 2622 472
rect 2522 357 2535 403
rect 2581 357 2622 403
rect 2522 288 2622 357
rect 2390 267 2438 288
rect 2318 228 2438 267
rect 2502 228 2622 288
rect 131 24 251 68
rect 299 24 419 68
rect 577 24 697 68
rect 759 24 879 68
rect 1071 24 1191 68
rect 1275 24 1395 68
rect 1499 24 1619 68
rect 1683 24 1803 68
rect 1910 24 2030 68
rect 2094 24 2214 68
rect 2318 24 2438 68
rect 2502 24 2622 68
<< polycontact >>
rect 155 393 201 439
rect 764 393 810 439
rect 312 261 358 307
rect 614 268 660 314
rect 1308 393 1354 439
rect 1132 265 1178 311
rect 1696 347 1742 393
rect 1951 393 1997 439
rect 2144 267 2190 313
rect 2344 267 2390 313
rect 2535 357 2581 403
<< metal1 >>
rect 0 724 2800 844
rect 45 665 113 724
rect 45 525 56 665
rect 102 525 113 665
rect 45 506 113 525
rect 249 665 317 676
rect 249 525 260 665
rect 306 552 317 665
rect 464 665 510 724
rect 464 608 510 619
rect 657 665 725 676
rect 657 552 668 665
rect 306 525 668 552
rect 714 552 725 665
rect 872 665 918 724
rect 1004 632 1016 678
rect 1062 632 1424 678
rect 1470 632 1832 678
rect 1878 632 2243 678
rect 2289 632 2651 678
rect 2697 632 2710 678
rect 872 608 918 619
rect 714 525 1220 552
rect 249 506 1220 525
rect 1266 506 1628 552
rect 1674 506 1685 552
rect 1810 488 2039 534
rect 2085 488 2447 534
rect 2493 488 2697 534
rect 131 393 155 439
rect 201 393 764 439
rect 810 393 831 439
rect 445 360 831 393
rect 914 393 1308 439
rect 1354 393 1365 439
rect 914 357 1365 393
rect 1474 393 1742 430
rect 914 354 1092 357
rect 1474 347 1696 393
rect 130 314 358 318
rect 130 307 614 314
rect 130 261 312 307
rect 358 268 614 307
rect 660 268 697 314
rect 1474 311 1742 347
rect 1121 265 1132 311
rect 1178 265 1742 311
rect 130 242 358 261
rect 1810 219 1894 488
rect 1940 393 1951 439
rect 1997 403 2592 439
rect 1997 393 2535 403
rect 1940 392 2535 393
rect 2488 357 2535 392
rect 2581 357 2592 403
rect 1974 313 2401 326
rect 1974 267 2144 313
rect 2190 267 2344 313
rect 2390 267 2401 313
rect 1974 242 2401 267
rect 404 215 1894 219
rect 404 194 996 215
rect 45 148 56 194
rect 102 173 996 194
rect 102 148 450 173
rect 985 169 996 173
rect 1042 173 1832 215
rect 1042 169 1053 173
rect 1810 169 1832 173
rect 1878 169 1894 215
rect 1810 158 1894 169
rect 491 81 502 127
rect 548 81 559 127
rect 491 60 559 81
rect 1413 81 1424 127
rect 1470 81 1481 127
rect 1413 60 1481 81
rect 2232 81 2243 127
rect 2289 81 2300 127
rect 2488 110 2592 357
rect 2651 171 2697 488
rect 2651 114 2697 125
rect 2232 60 2300 81
rect 0 -60 2800 60
<< labels >>
flabel metal1 s 914 357 1365 439 0 FreeSans 400 0 0 0 B2
port 4 nsew default input
flabel metal1 s 1474 311 1742 430 0 FreeSans 400 0 0 0 B1
port 3 nsew default input
flabel metal1 s 1974 242 2401 326 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1940 392 2592 439 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1810 488 2697 534 0 FreeSans 400 0 0 0 ZN
port 7 nsew default output
flabel metal1 s 2232 60 2300 127 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 0 724 2800 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 130 314 358 318 0 FreeSans 400 0 0 0 C2
port 6 nsew default input
flabel metal1 s 131 393 831 439 0 FreeSans 400 0 0 0 C1
port 5 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 2488 110 2592 392 1 A1
port 1 nsew default input
rlabel metal1 s 1121 265 1742 311 1 B1
port 3 nsew default input
rlabel metal1 s 914 354 1092 357 1 B2
port 4 nsew default input
rlabel metal1 s 445 360 831 393 1 C1
port 5 nsew default input
rlabel metal1 s 130 268 697 314 1 C2
port 6 nsew default input
rlabel metal1 s 130 242 358 268 1 C2
port 6 nsew default input
rlabel metal1 s 2651 219 2697 488 1 ZN
port 7 nsew default output
rlabel metal1 s 1810 219 1894 488 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 194 2697 219 1 ZN
port 7 nsew default output
rlabel metal1 s 404 194 1894 219 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 173 2697 194 1 ZN
port 7 nsew default output
rlabel metal1 s 45 173 1894 194 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 169 2697 173 1 ZN
port 7 nsew default output
rlabel metal1 s 1810 169 1894 173 1 ZN
port 7 nsew default output
rlabel metal1 s 985 169 1053 173 1 ZN
port 7 nsew default output
rlabel metal1 s 45 169 450 173 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 158 2697 169 1 ZN
port 7 nsew default output
rlabel metal1 s 1810 158 1894 169 1 ZN
port 7 nsew default output
rlabel metal1 s 45 158 450 169 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 148 2697 158 1 ZN
port 7 nsew default output
rlabel metal1 s 45 148 450 158 1 ZN
port 7 nsew default output
rlabel metal1 s 2651 114 2697 148 1 ZN
port 7 nsew default output
rlabel metal1 s 872 608 918 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 464 608 510 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 45 608 113 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 45 506 113 608 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1413 60 1481 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 491 60 559 127 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2800 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2800 784
string GDS_END 1294366
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1288452
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
