magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -80 2472 80 2531
rect -80 2426 -23 2472
rect 23 2426 80 2472
rect -80 2308 80 2426
rect -80 2262 -23 2308
rect 23 2262 80 2308
rect -80 2145 80 2262
rect -80 2099 -23 2145
rect 23 2099 80 2145
rect -80 1982 80 2099
rect -80 1936 -23 1982
rect 23 1936 80 1982
rect -80 1819 80 1936
rect -80 1773 -23 1819
rect 23 1773 80 1819
rect -80 1656 80 1773
rect -80 1610 -23 1656
rect 23 1610 80 1656
rect -80 1492 80 1610
rect -80 1446 -23 1492
rect 23 1446 80 1492
rect -80 1329 80 1446
rect -80 1283 -23 1329
rect 23 1283 80 1329
rect -80 1166 80 1283
rect -80 1120 -23 1166
rect 23 1120 80 1166
rect -80 1003 80 1120
rect -80 957 -23 1003
rect 23 957 80 1003
rect -80 839 80 957
rect -80 793 -23 839
rect 23 793 80 839
rect -80 676 80 793
rect -80 630 -23 676
rect 23 630 80 676
rect -80 513 80 630
rect -80 467 -23 513
rect 23 467 80 513
rect -80 350 80 467
rect -80 304 -23 350
rect 23 304 80 350
rect -80 186 80 304
rect -80 140 -23 186
rect 23 140 80 186
rect -80 23 80 140
rect -80 -23 -23 23
rect 23 -23 80 23
rect -80 -140 80 -23
rect -80 -186 -23 -140
rect 23 -186 80 -140
rect -80 -304 80 -186
rect -80 -350 -23 -304
rect 23 -350 80 -304
rect -80 -467 80 -350
rect -80 -513 -23 -467
rect 23 -513 80 -467
rect -80 -630 80 -513
rect -80 -676 -23 -630
rect 23 -676 80 -630
rect -80 -793 80 -676
rect -80 -839 -23 -793
rect 23 -839 80 -793
rect -80 -957 80 -839
rect -80 -1003 -23 -957
rect 23 -1003 80 -957
rect -80 -1120 80 -1003
rect -80 -1166 -23 -1120
rect 23 -1166 80 -1120
rect -80 -1283 80 -1166
rect -80 -1329 -23 -1283
rect 23 -1329 80 -1283
rect -80 -1446 80 -1329
rect -80 -1492 -23 -1446
rect 23 -1492 80 -1446
rect -80 -1610 80 -1492
rect -80 -1656 -23 -1610
rect 23 -1656 80 -1610
rect -80 -1773 80 -1656
rect -80 -1819 -23 -1773
rect 23 -1819 80 -1773
rect -80 -1936 80 -1819
rect -80 -1982 -23 -1936
rect 23 -1982 80 -1936
rect -80 -2099 80 -1982
rect -80 -2145 -23 -2099
rect 23 -2145 80 -2099
rect -80 -2262 80 -2145
rect -80 -2308 -23 -2262
rect 23 -2308 80 -2262
rect -80 -2426 80 -2308
rect -80 -2472 -23 -2426
rect 23 -2472 80 -2426
rect -80 -2530 80 -2472
<< psubdiffcont >>
rect -23 2426 23 2472
rect -23 2262 23 2308
rect -23 2099 23 2145
rect -23 1936 23 1982
rect -23 1773 23 1819
rect -23 1610 23 1656
rect -23 1446 23 1492
rect -23 1283 23 1329
rect -23 1120 23 1166
rect -23 957 23 1003
rect -23 793 23 839
rect -23 630 23 676
rect -23 467 23 513
rect -23 304 23 350
rect -23 140 23 186
rect -23 -23 23 23
rect -23 -186 23 -140
rect -23 -350 23 -304
rect -23 -513 23 -467
rect -23 -676 23 -630
rect -23 -839 23 -793
rect -23 -1003 23 -957
rect -23 -1166 23 -1120
rect -23 -1329 23 -1283
rect -23 -1492 23 -1446
rect -23 -1656 23 -1610
rect -23 -1819 23 -1773
rect -23 -1982 23 -1936
rect -23 -2145 23 -2099
rect -23 -2308 23 -2262
rect -23 -2472 23 -2426
<< metal1 >>
rect -71 2472 71 2522
rect -71 2426 -23 2472
rect 23 2426 71 2472
rect -71 2308 71 2426
rect -71 2262 -23 2308
rect 23 2262 71 2308
rect -71 2145 71 2262
rect -71 2099 -23 2145
rect 23 2099 71 2145
rect -71 1982 71 2099
rect -71 1936 -23 1982
rect 23 1936 71 1982
rect -71 1819 71 1936
rect -71 1773 -23 1819
rect 23 1773 71 1819
rect -71 1656 71 1773
rect -71 1610 -23 1656
rect 23 1610 71 1656
rect -71 1492 71 1610
rect -71 1446 -23 1492
rect 23 1446 71 1492
rect -71 1329 71 1446
rect -71 1283 -23 1329
rect 23 1283 71 1329
rect -71 1166 71 1283
rect -71 1120 -23 1166
rect 23 1120 71 1166
rect -71 1003 71 1120
rect -71 957 -23 1003
rect 23 957 71 1003
rect -71 839 71 957
rect -71 793 -23 839
rect 23 793 71 839
rect -71 676 71 793
rect -71 630 -23 676
rect 23 630 71 676
rect -71 513 71 630
rect -71 467 -23 513
rect 23 467 71 513
rect -71 350 71 467
rect -71 304 -23 350
rect 23 304 71 350
rect -71 186 71 304
rect -71 140 -23 186
rect 23 140 71 186
rect -71 23 71 140
rect -71 -23 -23 23
rect 23 -23 71 23
rect -71 -140 71 -23
rect -71 -186 -23 -140
rect 23 -186 71 -140
rect -71 -304 71 -186
rect -71 -350 -23 -304
rect 23 -350 71 -304
rect -71 -467 71 -350
rect -71 -513 -23 -467
rect 23 -513 71 -467
rect -71 -630 71 -513
rect -71 -676 -23 -630
rect 23 -676 71 -630
rect -71 -793 71 -676
rect -71 -839 -23 -793
rect 23 -839 71 -793
rect -71 -957 71 -839
rect -71 -1003 -23 -957
rect 23 -1003 71 -957
rect -71 -1120 71 -1003
rect -71 -1166 -23 -1120
rect 23 -1166 71 -1120
rect -71 -1283 71 -1166
rect -71 -1329 -23 -1283
rect 23 -1329 71 -1283
rect -71 -1446 71 -1329
rect -71 -1492 -23 -1446
rect 23 -1492 71 -1446
rect -71 -1610 71 -1492
rect -71 -1656 -23 -1610
rect 23 -1656 71 -1610
rect -71 -1773 71 -1656
rect -71 -1819 -23 -1773
rect 23 -1819 71 -1773
rect -71 -1936 71 -1819
rect -71 -1982 -23 -1936
rect 23 -1982 71 -1936
rect -71 -2099 71 -1982
rect -71 -2145 -23 -2099
rect 23 -2145 71 -2099
rect -71 -2262 71 -2145
rect -71 -2308 -23 -2262
rect 23 -2308 71 -2262
rect -71 -2426 71 -2308
rect -71 -2472 -23 -2426
rect 23 -2472 71 -2426
rect -71 -2522 71 -2472
<< properties >>
string GDS_END 311110
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 308930
<< end >>
