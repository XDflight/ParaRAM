magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 124 116 244 300
rect 348 116 468 300
rect 572 116 692 300
rect 796 116 916 300
<< mvpmos >>
rect 134 573 234 939
rect 358 573 458 939
rect 572 573 672 939
rect 806 573 906 939
<< mvndiff >>
rect 36 269 124 300
rect 36 129 49 269
rect 95 129 124 269
rect 36 116 124 129
rect 244 287 348 300
rect 244 147 273 287
rect 319 147 348 287
rect 244 116 348 147
rect 468 175 572 300
rect 468 129 497 175
rect 543 129 572 175
rect 468 116 572 129
rect 692 287 796 300
rect 692 147 721 287
rect 767 147 796 287
rect 692 116 796 147
rect 916 269 1004 300
rect 916 129 945 269
rect 991 129 1004 269
rect 916 116 1004 129
<< mvpdiff >>
rect 46 861 134 939
rect 46 721 59 861
rect 105 721 134 861
rect 46 573 134 721
rect 234 573 358 939
rect 458 861 572 939
rect 458 721 497 861
rect 543 721 572 861
rect 458 573 572 721
rect 672 573 806 939
rect 906 861 994 939
rect 906 721 935 861
rect 981 721 994 861
rect 906 573 994 721
<< mvndiffc >>
rect 49 129 95 269
rect 273 147 319 287
rect 497 129 543 175
rect 721 147 767 287
rect 945 129 991 269
<< mvpdiffc >>
rect 59 721 105 861
rect 497 721 543 861
rect 935 721 981 861
<< polysilicon >>
rect 134 939 234 983
rect 358 939 458 983
rect 572 939 672 983
rect 806 939 906 983
rect 134 500 234 573
rect 134 454 175 500
rect 221 454 234 500
rect 134 344 234 454
rect 358 513 458 573
rect 572 513 672 573
rect 806 513 906 573
rect 358 500 672 513
rect 358 454 371 500
rect 417 454 672 500
rect 358 441 672 454
rect 720 500 906 513
rect 720 454 733 500
rect 779 454 906 500
rect 720 441 906 454
rect 358 344 468 441
rect 124 300 244 344
rect 348 300 468 344
rect 572 344 672 441
rect 796 344 906 441
rect 572 300 692 344
rect 796 300 916 344
rect 124 72 244 116
rect 348 72 468 116
rect 572 72 692 116
rect 796 72 916 116
<< polycontact >>
rect 175 454 221 500
rect 371 454 417 500
rect 733 454 779 500
<< metal1 >>
rect 0 918 1120 1098
rect 59 861 105 918
rect 59 710 105 721
rect 497 861 543 872
rect 935 861 981 918
rect 543 721 882 756
rect 497 710 882 721
rect 935 710 981 721
rect 175 588 790 634
rect 175 500 221 588
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 702 500 790 588
rect 702 454 733 500
rect 779 454 790 500
rect 175 443 221 454
rect 702 354 754 454
rect 836 344 882 710
rect 814 298 882 344
rect 273 287 882 298
rect 49 269 95 280
rect 319 232 721 287
rect 273 136 319 147
rect 497 175 543 186
rect 49 90 95 129
rect 767 242 882 287
rect 945 269 991 280
rect 721 136 767 147
rect 497 90 543 129
rect 945 90 991 129
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 175 588 790 634 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 945 186 991 280 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 497 756 543 872 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 702 454 790 588 1 A2
port 2 nsew default input
rlabel metal1 s 175 454 221 588 1 A2
port 2 nsew default input
rlabel metal1 s 702 443 754 454 1 A2
port 2 nsew default input
rlabel metal1 s 175 443 221 454 1 A2
port 2 nsew default input
rlabel metal1 s 702 354 754 443 1 A2
port 2 nsew default input
rlabel metal1 s 497 710 882 756 1 ZN
port 3 nsew default output
rlabel metal1 s 836 344 882 710 1 ZN
port 3 nsew default output
rlabel metal1 s 814 298 882 344 1 ZN
port 3 nsew default output
rlabel metal1 s 273 242 882 298 1 ZN
port 3 nsew default output
rlabel metal1 s 273 232 767 242 1 ZN
port 3 nsew default output
rlabel metal1 s 721 136 767 232 1 ZN
port 3 nsew default output
rlabel metal1 s 273 136 319 232 1 ZN
port 3 nsew default output
rlabel metal1 s 935 710 981 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 59 710 105 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 49 186 95 280 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 186 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 497 90 543 186 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 186 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 78802
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 75422
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
