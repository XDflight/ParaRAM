magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 396 5574 870
rect -86 352 1977 396
rect 3404 352 5574 396
<< pwell >>
rect 1977 352 3404 396
rect -86 -86 5574 352
<< mvnmos >>
rect 124 151 244 232
rect 348 151 468 232
rect 740 156 860 232
rect 964 156 1084 232
rect 1188 156 1308 232
rect 1356 156 1476 232
rect 1888 156 2008 232
rect 2424 204 2544 276
rect 2634 204 2754 276
rect 2858 204 2978 276
rect 3082 204 3202 276
rect 3643 156 3763 228
rect 3811 156 3931 228
rect 4035 156 4155 228
rect 4203 156 4323 228
rect 4571 69 4691 232
rect 4795 69 4915 232
rect 5019 69 5139 232
rect 5243 69 5363 232
<< mvpmos >>
rect 144 487 244 660
rect 348 487 448 660
rect 740 504 840 586
rect 944 504 1044 586
rect 1148 504 1248 586
rect 1356 504 1456 586
rect 1984 516 2084 677
rect 2444 516 2544 677
rect 2809 516 2909 628
rect 3013 516 3113 628
rect 3217 516 3317 628
rect 3627 472 3727 647
rect 3831 472 3931 647
rect 4035 472 4135 647
rect 4239 472 4339 647
rect 4591 472 4691 715
rect 4795 472 4895 715
rect 4999 472 5099 715
rect 5203 472 5303 715
<< mvndiff >>
rect 2161 232 2424 276
rect 36 219 124 232
rect 36 173 49 219
rect 95 173 124 219
rect 36 151 124 173
rect 244 210 348 232
rect 244 164 273 210
rect 319 164 348 210
rect 244 151 348 164
rect 468 219 556 232
rect 468 173 497 219
rect 543 173 556 219
rect 468 151 556 173
rect 652 215 740 232
rect 652 169 665 215
rect 711 169 740 215
rect 652 156 740 169
rect 860 215 964 232
rect 860 169 889 215
rect 935 169 964 215
rect 860 156 964 169
rect 1084 215 1188 232
rect 1084 169 1113 215
rect 1159 169 1188 215
rect 1084 156 1188 169
rect 1308 156 1356 232
rect 1476 156 1888 232
rect 2008 204 2424 232
rect 2544 204 2634 276
rect 2754 263 2858 276
rect 2754 217 2783 263
rect 2829 217 2858 263
rect 2754 204 2858 217
rect 2978 263 3082 276
rect 2978 217 3007 263
rect 3053 217 3082 263
rect 2978 204 3082 217
rect 3202 263 3293 276
rect 3202 217 3234 263
rect 3280 217 3293 263
rect 3202 204 3293 217
rect 2008 183 2364 204
rect 2008 156 2127 183
rect 2114 137 2127 156
rect 2173 152 2364 183
rect 2173 137 2186 152
rect 2114 124 2186 137
rect 3555 215 3643 228
rect 3555 169 3568 215
rect 3614 169 3643 215
rect 3555 156 3643 169
rect 3763 156 3811 228
rect 3931 215 4035 228
rect 3931 169 3960 215
rect 4006 169 4035 215
rect 3931 156 4035 169
rect 4155 156 4203 228
rect 4323 215 4411 228
rect 4323 169 4352 215
rect 4398 169 4411 215
rect 4323 156 4411 169
rect 4483 142 4571 232
rect 4483 96 4496 142
rect 4542 96 4571 142
rect 4483 69 4571 96
rect 4691 167 4795 232
rect 4691 121 4720 167
rect 4766 121 4795 167
rect 4691 69 4795 121
rect 4915 142 5019 232
rect 4915 96 4944 142
rect 4990 96 5019 142
rect 4915 69 5019 96
rect 5139 167 5243 232
rect 5139 121 5168 167
rect 5214 121 5243 167
rect 5139 69 5243 121
rect 5363 142 5451 232
rect 5363 96 5392 142
rect 5438 96 5451 142
rect 5363 69 5451 96
<< mvpdiff >>
rect 56 647 144 660
rect 56 507 69 647
rect 115 507 144 647
rect 56 487 144 507
rect 244 647 348 660
rect 244 601 273 647
rect 319 601 348 647
rect 244 487 348 601
rect 448 647 536 660
rect 448 507 477 647
rect 523 507 536 647
rect 448 487 536 507
rect 608 646 680 659
rect 608 600 621 646
rect 667 600 680 646
rect 608 586 680 600
rect 1516 679 1588 692
rect 1516 633 1529 679
rect 1575 677 1588 679
rect 1575 633 1984 677
rect 1516 586 1984 633
rect 608 504 740 586
rect 840 566 944 586
rect 840 520 869 566
rect 915 520 944 566
rect 840 504 944 520
rect 1044 566 1148 586
rect 1044 520 1073 566
rect 1119 520 1148 566
rect 1044 504 1148 520
rect 1248 563 1356 586
rect 1248 517 1281 563
rect 1327 517 1356 563
rect 1248 504 1356 517
rect 1456 516 1984 586
rect 2084 575 2172 677
rect 2084 529 2113 575
rect 2159 529 2172 575
rect 2084 516 2172 529
rect 2356 575 2444 677
rect 2356 529 2369 575
rect 2415 529 2444 575
rect 2356 516 2444 529
rect 2544 664 2749 677
rect 2544 618 2690 664
rect 2736 628 2749 664
rect 4503 665 4591 715
rect 3539 634 3627 647
rect 2736 618 2809 628
rect 2544 516 2809 618
rect 2909 575 3013 628
rect 2909 529 2938 575
rect 2984 529 3013 575
rect 2909 516 3013 529
rect 3113 579 3217 628
rect 3113 533 3142 579
rect 3188 533 3217 579
rect 3113 516 3217 533
rect 3317 579 3405 628
rect 3317 533 3346 579
rect 3392 533 3405 579
rect 3317 516 3405 533
rect 3539 588 3552 634
rect 3598 588 3627 634
rect 1456 504 1700 516
rect 3539 472 3627 588
rect 3727 560 3831 647
rect 3727 514 3756 560
rect 3802 514 3831 560
rect 3727 472 3831 514
rect 3931 634 4035 647
rect 3931 588 3960 634
rect 4006 588 4035 634
rect 3931 472 4035 588
rect 4135 560 4239 647
rect 4135 514 4164 560
rect 4210 514 4239 560
rect 4135 472 4239 514
rect 4339 634 4427 647
rect 4339 494 4368 634
rect 4414 494 4427 634
rect 4339 472 4427 494
rect 4503 525 4516 665
rect 4562 525 4591 665
rect 4503 472 4591 525
rect 4691 665 4795 715
rect 4691 525 4720 665
rect 4766 525 4795 665
rect 4691 472 4795 525
rect 4895 665 4999 715
rect 4895 525 4924 665
rect 4970 525 4999 665
rect 4895 472 4999 525
rect 5099 665 5203 715
rect 5099 525 5128 665
rect 5174 525 5203 665
rect 5099 472 5203 525
rect 5303 665 5391 715
rect 5303 525 5332 665
rect 5378 525 5391 665
rect 5303 472 5391 525
<< mvndiffc >>
rect 49 173 95 219
rect 273 164 319 210
rect 497 173 543 219
rect 665 169 711 215
rect 889 169 935 215
rect 1113 169 1159 215
rect 2783 217 2829 263
rect 3007 217 3053 263
rect 3234 217 3280 263
rect 2127 137 2173 183
rect 3568 169 3614 215
rect 3960 169 4006 215
rect 4352 169 4398 215
rect 4496 96 4542 142
rect 4720 121 4766 167
rect 4944 96 4990 142
rect 5168 121 5214 167
rect 5392 96 5438 142
<< mvpdiffc >>
rect 69 507 115 647
rect 273 601 319 647
rect 477 507 523 647
rect 621 600 667 646
rect 1529 633 1575 679
rect 869 520 915 566
rect 1073 520 1119 566
rect 1281 517 1327 563
rect 2113 529 2159 575
rect 2369 529 2415 575
rect 2690 618 2736 664
rect 2938 529 2984 575
rect 3142 533 3188 579
rect 3346 533 3392 579
rect 3552 588 3598 634
rect 3756 514 3802 560
rect 3960 588 4006 634
rect 4164 514 4210 560
rect 4368 494 4414 634
rect 4516 525 4562 665
rect 4720 525 4766 665
rect 4924 525 4970 665
rect 5128 525 5174 665
rect 5332 525 5378 665
<< polysilicon >>
rect 348 720 1044 760
rect 144 660 244 704
rect 348 660 448 720
rect 740 586 840 630
rect 944 586 1044 720
rect 1148 667 1248 680
rect 1148 621 1161 667
rect 1207 621 1248 667
rect 1984 677 2084 721
rect 2444 677 2544 721
rect 2809 720 3727 760
rect 1148 586 1248 621
rect 1356 586 1456 630
rect 2809 628 2909 720
rect 3013 628 3113 672
rect 3217 628 3317 672
rect 3627 647 3727 720
rect 4591 715 4691 760
rect 4795 715 4895 760
rect 4999 715 5099 760
rect 5203 715 5303 760
rect 3831 647 3931 691
rect 4035 647 4135 691
rect 4239 647 4339 691
rect 144 418 244 487
rect 144 372 157 418
rect 203 372 244 418
rect 144 276 244 372
rect 124 232 244 276
rect 348 323 448 487
rect 348 277 365 323
rect 411 277 448 323
rect 348 276 448 277
rect 740 415 840 504
rect 944 460 1044 504
rect 740 369 753 415
rect 799 369 840 415
rect 1148 428 1248 504
rect 1356 444 1456 504
rect 1148 412 1188 428
rect 740 292 840 369
rect 964 372 1188 412
rect 348 232 468 276
rect 740 232 860 292
rect 964 232 1084 372
rect 1225 311 1308 324
rect 1225 292 1238 311
rect 1188 265 1238 292
rect 1284 265 1308 311
rect 1188 232 1308 265
rect 1356 311 1476 444
rect 1984 427 2084 516
rect 2444 456 2544 516
rect 1356 265 1417 311
rect 1463 265 1476 311
rect 1356 232 1476 265
rect 1888 387 2084 427
rect 1888 232 2008 387
rect 2424 355 2544 456
rect 2809 444 2909 516
rect 2424 309 2437 355
rect 2483 309 2544 355
rect 2424 276 2544 309
rect 2634 404 2909 444
rect 3013 471 3113 516
rect 3013 425 3050 471
rect 3096 444 3113 471
rect 3217 460 3317 516
rect 3277 444 3317 460
rect 3096 425 3122 444
rect 2634 276 2754 404
rect 3013 392 3122 425
rect 3277 404 3425 444
rect 3627 418 3727 472
rect 3082 344 3122 392
rect 2858 276 2978 344
rect 3082 276 3202 344
rect 124 107 244 151
rect 348 64 468 151
rect 740 112 860 156
rect 964 112 1084 156
rect 1188 64 1308 156
rect 1356 112 1476 156
rect 348 24 1308 64
rect 1888 64 2008 156
rect 2424 152 2544 204
rect 2634 152 2754 204
rect 2858 171 2978 204
rect 2858 125 2897 171
rect 2943 125 2978 171
rect 3082 152 3202 204
rect 3353 171 3425 404
rect 3643 415 3727 418
rect 3643 275 3656 415
rect 3702 275 3727 415
rect 3643 272 3727 275
rect 3831 308 3931 472
rect 3831 272 3872 308
rect 3643 228 3763 272
rect 3811 262 3872 272
rect 3918 262 3931 308
rect 3811 228 3931 262
rect 4035 415 4135 472
rect 4035 369 4048 415
rect 4094 369 4135 415
rect 4035 272 4135 369
rect 4239 439 4339 472
rect 4239 393 4276 439
rect 4322 393 4339 439
rect 4239 380 4339 393
rect 4239 272 4323 380
rect 4591 357 4691 472
rect 4795 357 4895 472
rect 4999 357 5099 472
rect 5203 357 5303 472
rect 4591 353 5303 357
rect 4591 307 4604 353
rect 4650 311 4823 353
rect 4650 307 4691 311
rect 4591 276 4691 307
rect 4035 228 4155 272
rect 4203 228 4323 272
rect 4571 232 4691 276
rect 4795 307 4823 311
rect 4869 311 5032 353
rect 4869 307 4915 311
rect 4795 232 4915 307
rect 5019 307 5032 311
rect 5078 311 5303 353
rect 5078 307 5139 311
rect 5019 232 5139 307
rect 5243 276 5303 311
rect 5243 232 5363 276
rect 2858 112 2978 125
rect 3353 125 3366 171
rect 3412 125 3425 171
rect 3353 112 3425 125
rect 3643 112 3763 156
rect 3811 112 3931 156
rect 4035 64 4155 156
rect 4203 112 4323 156
rect 1888 24 4155 64
rect 4571 24 4691 69
rect 4795 24 4915 69
rect 5019 24 5139 69
rect 5243 24 5363 69
<< polycontact >>
rect 1161 621 1207 667
rect 157 372 203 418
rect 365 277 411 323
rect 753 369 799 415
rect 1238 265 1284 311
rect 1417 265 1463 311
rect 2437 309 2483 355
rect 3050 425 3096 471
rect 2897 125 2943 171
rect 3656 275 3702 415
rect 3872 262 3918 308
rect 4048 369 4094 415
rect 4276 393 4322 439
rect 4604 307 4650 353
rect 4823 307 4869 353
rect 5032 307 5078 353
rect 3366 125 3412 171
<< metal1 >>
rect 0 724 5488 844
rect 69 647 115 660
rect 262 647 330 724
rect 262 601 273 647
rect 319 601 330 647
rect 477 647 523 660
rect 115 507 411 534
rect 69 487 411 507
rect 56 418 318 430
rect 56 372 157 418
rect 203 372 318 418
rect 56 354 318 372
rect 365 323 411 487
rect 49 277 365 302
rect 49 256 411 277
rect 610 646 678 724
rect 1517 679 1586 724
rect 610 600 621 646
rect 667 600 678 646
rect 757 621 1161 667
rect 1207 621 1419 667
rect 1517 633 1529 679
rect 1575 633 1586 679
rect 757 554 803 621
rect 1373 587 1419 621
rect 1656 632 2644 678
rect 1656 587 1702 632
rect 523 508 803 554
rect 858 520 869 566
rect 915 520 946 566
rect 49 219 95 256
rect 477 230 523 507
rect 578 415 810 430
rect 578 369 753 415
rect 799 369 810 415
rect 578 354 810 369
rect 477 219 543 230
rect 49 162 95 173
rect 262 164 273 210
rect 319 164 330 210
rect 262 60 330 164
rect 477 173 497 219
rect 858 215 946 520
rect 1062 520 1073 566
rect 1119 520 1130 566
rect 1062 403 1130 520
rect 1281 563 1327 574
rect 1373 541 1702 587
rect 2102 563 2113 575
rect 1281 495 1327 517
rect 1748 529 2113 563
rect 2159 529 2170 575
rect 2358 529 2369 575
rect 2415 529 2552 575
rect 1748 517 2170 529
rect 1748 495 1794 517
rect 1281 449 1794 495
rect 2506 469 2552 529
rect 2598 561 2644 632
rect 2690 664 2736 724
rect 2690 607 2736 618
rect 2835 632 3096 678
rect 2835 561 2881 632
rect 2598 515 2881 561
rect 2927 529 2938 575
rect 2984 529 2995 575
rect 2927 469 2995 529
rect 1840 414 2460 460
rect 2506 425 2995 469
rect 3050 471 3096 632
rect 2506 423 2950 425
rect 1840 403 1886 414
rect 1062 357 1886 403
rect 477 162 543 173
rect 654 169 665 215
rect 711 169 722 215
rect 858 169 889 215
rect 935 169 946 215
rect 1113 215 1159 357
rect 1932 321 2368 367
rect 1932 311 1978 321
rect 654 60 722 169
rect 1113 158 1159 169
rect 1227 265 1238 311
rect 1284 265 1295 311
rect 1406 265 1417 311
rect 1463 265 1978 311
rect 1227 204 1295 265
rect 2024 229 2276 275
rect 2024 204 2070 229
rect 1227 158 2070 204
rect 2116 137 2127 183
rect 2173 137 2184 183
rect 2116 60 2184 137
rect 2230 152 2276 229
rect 2322 263 2368 321
rect 2414 355 2460 414
rect 2414 309 2437 355
rect 2483 309 2494 355
rect 2893 263 2950 423
rect 3050 414 3096 425
rect 3142 632 3495 678
rect 3142 579 3188 632
rect 3142 263 3188 533
rect 3335 533 3346 579
rect 3392 533 3403 579
rect 3335 274 3403 533
rect 3449 542 3495 632
rect 3541 634 3609 724
rect 3541 588 3552 634
rect 3598 588 3609 634
rect 3655 617 3894 664
rect 3655 542 3701 617
rect 3449 495 3701 542
rect 3756 560 3802 571
rect 3490 415 3708 430
rect 3490 354 3656 415
rect 2322 217 2783 263
rect 2829 217 2950 263
rect 2996 217 3007 263
rect 3053 217 3188 263
rect 3234 263 3403 274
rect 3645 275 3656 354
rect 3702 275 3708 415
rect 3645 264 3708 275
rect 3280 217 3592 263
rect 3234 206 3291 217
rect 3535 215 3592 217
rect 3756 215 3802 514
rect 3848 542 3894 617
rect 3949 634 4017 724
rect 3949 588 3960 634
rect 4006 588 4017 634
rect 4063 617 4322 664
rect 4063 542 4109 617
rect 3848 496 4109 542
rect 4164 560 4230 571
rect 4210 514 4230 560
rect 4164 503 4230 514
rect 3876 415 4126 430
rect 3876 369 4048 415
rect 4094 369 4126 415
rect 3876 354 4126 369
rect 4184 312 4230 503
rect 4276 439 4322 617
rect 4368 634 4414 724
rect 4516 665 4562 724
rect 4516 514 4562 525
rect 4709 665 4777 676
rect 4709 525 4720 665
rect 4766 525 4777 665
rect 4368 483 4414 494
rect 4709 466 4777 525
rect 4924 665 4970 724
rect 4924 514 4970 525
rect 5117 665 5246 676
rect 5117 525 5128 665
rect 5174 525 5246 665
rect 5117 466 5246 525
rect 5332 665 5378 724
rect 5332 514 5378 525
rect 4709 420 5246 466
rect 4276 382 4322 393
rect 4593 353 5078 364
rect 4593 312 4604 353
rect 4184 308 4604 312
rect 3861 262 3872 308
rect 3918 307 4604 308
rect 4650 307 4823 353
rect 4869 307 5032 353
rect 3918 295 5078 307
rect 3918 266 4661 295
rect 3918 262 4398 266
rect 4352 215 4398 262
rect 5170 234 5246 420
rect 2886 152 2897 171
rect 2230 125 2897 152
rect 2943 152 2954 171
rect 3355 152 3366 171
rect 2943 125 3366 152
rect 3412 125 3423 171
rect 3535 169 3568 215
rect 3614 169 3802 215
rect 3535 158 3802 169
rect 3949 169 3960 215
rect 4006 169 4017 215
rect 2230 106 3423 125
rect 3949 60 4017 169
rect 4352 158 4398 169
rect 4720 188 5246 234
rect 4720 167 4766 188
rect 4496 142 4542 153
rect 5168 167 5246 188
rect 4720 110 4766 121
rect 4496 60 4542 96
rect 4933 96 4944 142
rect 4990 96 5001 142
rect 5214 121 5246 167
rect 5168 110 5246 121
rect 5392 142 5438 153
rect 4933 60 5001 96
rect 5392 60 5438 96
rect 0 -60 5488 60
<< labels >>
flabel metal1 s 578 354 810 430 0 FreeSans 600 0 0 0 D
port 1 nsew default input
flabel metal1 s 5117 466 5246 676 0 FreeSans 600 0 0 0 Q
port 5 nsew default output
flabel metal1 s 3876 354 4126 430 0 FreeSans 600 0 0 0 RN
port 2 nsew default input
flabel metal1 s 3490 354 3708 430 0 FreeSans 600 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 0 724 5488 844 0 FreeSans 600 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3949 210 4017 215 0 FreeSans 600 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 56 354 318 430 0 FreeSans 600 0 0 0 CLKN
port 4 nsew clock input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3645 264 3708 354 1 SETN
port 3 nsew default input
rlabel metal1 s 4709 466 4777 676 1 Q
port 5 nsew default output
rlabel metal1 s 4709 420 5246 466 1 Q
port 5 nsew default output
rlabel metal1 s 5170 234 5246 420 1 Q
port 5 nsew default output
rlabel metal1 s 4720 188 5246 234 1 Q
port 5 nsew default output
rlabel metal1 s 5168 110 5246 188 1 Q
port 5 nsew default output
rlabel metal1 s 4720 110 4766 188 1 Q
port 5 nsew default output
rlabel metal1 s 5332 633 5378 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 633 4970 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 633 4562 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 633 4414 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 633 4017 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 633 3609 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2690 633 2736 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1517 633 1586 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 633 678 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 633 330 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 607 5378 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 607 4970 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 607 4562 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 607 4414 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 607 4017 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 607 3609 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2690 607 2736 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 607 678 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 607 330 633 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 601 5378 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 601 4970 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 601 4562 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 601 4414 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 601 4017 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 601 3609 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 601 678 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 262 601 330 607 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 600 5378 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 600 4970 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 600 4562 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 600 4414 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 600 4017 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 600 3609 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 610 600 678 601 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 588 5378 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 588 4970 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 588 4562 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 588 4414 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3949 588 4017 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3541 588 3609 600 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 5332 514 5378 588 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4924 514 4970 588 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4516 514 4562 588 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 514 4414 588 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4368 483 4414 514 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 654 210 722 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 183 4017 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 183 722 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 183 330 210 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 153 4017 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 153 2184 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 153 722 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 153 330 183 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5392 142 5438 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4496 142 4542 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 142 4017 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 142 2184 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 142 722 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 142 330 153 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 5392 60 5438 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4933 60 5001 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4496 60 4542 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3949 60 4017 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2116 60 2184 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 654 60 722 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 142 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5488 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5488 784
string GDS_END 922820
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 911874
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
