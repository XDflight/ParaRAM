magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 456 3558 1094
rect -86 453 86 456
rect 3386 453 3558 456
<< pwell >>
rect 949 453 1291 456
rect -86 -86 3558 453
<< mvnmos >>
rect 124 156 244 288
rect 348 156 468 288
rect 572 156 692 288
rect 796 156 916 288
rect 1056 156 1176 336
rect 1426 169 1546 301
rect 1650 169 1770 301
rect 2018 201 2138 333
rect 2242 201 2362 333
rect 2466 201 2586 333
rect 2690 201 2810 333
rect 2914 201 3034 333
rect 3138 201 3258 333
<< mvpmos >>
rect 134 669 234 852
rect 404 669 504 852
rect 608 669 708 852
rect 816 669 916 852
rect 1056 576 1156 852
rect 1436 669 1536 852
rect 1640 669 1740 852
rect 2058 669 2158 852
rect 2262 669 2362 852
rect 2466 669 2566 852
rect 2670 669 2770 852
rect 2874 669 2974 852
rect 3078 669 3178 852
<< mvndiff >>
rect 976 288 1056 336
rect 36 275 124 288
rect 36 229 49 275
rect 95 229 124 275
rect 36 156 124 229
rect 244 275 348 288
rect 244 229 273 275
rect 319 229 348 275
rect 244 156 348 229
rect 468 275 572 288
rect 468 229 497 275
rect 543 229 572 275
rect 468 156 572 229
rect 692 275 796 288
rect 692 229 721 275
rect 767 229 796 275
rect 692 156 796 229
rect 916 275 1056 288
rect 916 229 945 275
rect 991 229 1056 275
rect 916 156 1056 229
rect 1176 299 1264 336
rect 1176 253 1205 299
rect 1251 253 1264 299
rect 1176 156 1264 253
rect 1338 288 1426 301
rect 1338 242 1351 288
rect 1397 242 1426 288
rect 1338 169 1426 242
rect 1546 258 1650 301
rect 1546 212 1575 258
rect 1621 212 1650 258
rect 1546 169 1650 212
rect 1770 275 1858 301
rect 1770 229 1799 275
rect 1845 229 1858 275
rect 1770 169 1858 229
rect 1930 275 2018 333
rect 1930 229 1943 275
rect 1989 229 2018 275
rect 1930 201 2018 229
rect 2138 275 2242 333
rect 2138 229 2167 275
rect 2213 229 2242 275
rect 2138 201 2242 229
rect 2362 275 2466 333
rect 2362 229 2391 275
rect 2437 229 2466 275
rect 2362 201 2466 229
rect 2586 275 2690 333
rect 2586 229 2615 275
rect 2661 229 2690 275
rect 2586 201 2690 229
rect 2810 275 2914 333
rect 2810 229 2839 275
rect 2885 229 2914 275
rect 2810 201 2914 229
rect 3034 275 3138 333
rect 3034 229 3063 275
rect 3109 229 3138 275
rect 3034 201 3138 229
rect 3258 275 3346 333
rect 3258 229 3287 275
rect 3333 229 3346 275
rect 3258 201 3346 229
<< mvpdiff >>
rect 46 839 134 852
rect 46 699 59 839
rect 105 699 134 839
rect 46 669 134 699
rect 234 823 404 852
rect 234 683 273 823
rect 319 683 404 823
rect 234 669 404 683
rect 504 823 608 852
rect 504 683 533 823
rect 579 683 608 823
rect 504 669 608 683
rect 708 728 816 852
rect 708 682 737 728
rect 783 682 816 728
rect 708 669 816 682
rect 916 830 1056 852
rect 916 784 945 830
rect 991 784 1056 830
rect 916 669 1056 784
rect 976 576 1056 669
rect 1156 635 1244 852
rect 1348 823 1436 852
rect 1348 683 1361 823
rect 1407 683 1436 823
rect 1348 669 1436 683
rect 1536 823 1640 852
rect 1536 683 1565 823
rect 1611 683 1640 823
rect 1536 669 1640 683
rect 1740 836 1828 852
rect 1740 696 1769 836
rect 1815 696 1828 836
rect 1740 669 1828 696
rect 1970 728 2058 852
rect 1970 682 1983 728
rect 2029 682 2058 728
rect 1970 669 2058 682
rect 2158 839 2262 852
rect 2158 699 2187 839
rect 2233 699 2262 839
rect 2158 669 2262 699
rect 2362 728 2466 852
rect 2362 682 2391 728
rect 2437 682 2466 728
rect 2362 669 2466 682
rect 2566 823 2670 852
rect 2566 683 2595 823
rect 2641 683 2670 823
rect 2566 669 2670 683
rect 2770 839 2874 852
rect 2770 699 2799 839
rect 2845 699 2874 839
rect 2770 669 2874 699
rect 2974 839 3078 852
rect 2974 699 3003 839
rect 3049 699 3078 839
rect 2974 669 3078 699
rect 3178 823 3266 852
rect 3178 683 3207 823
rect 3253 683 3266 823
rect 3178 669 3266 683
rect 1156 589 1185 635
rect 1231 589 1244 635
rect 1156 576 1244 589
<< mvndiffc >>
rect 49 229 95 275
rect 273 229 319 275
rect 497 229 543 275
rect 721 229 767 275
rect 945 229 991 275
rect 1205 253 1251 299
rect 1351 242 1397 288
rect 1575 212 1621 258
rect 1799 229 1845 275
rect 1943 229 1989 275
rect 2167 229 2213 275
rect 2391 229 2437 275
rect 2615 229 2661 275
rect 2839 229 2885 275
rect 3063 229 3109 275
rect 3287 229 3333 275
<< mvpdiffc >>
rect 59 699 105 839
rect 273 683 319 823
rect 533 683 579 823
rect 737 682 783 728
rect 945 784 991 830
rect 1361 683 1407 823
rect 1565 683 1611 823
rect 1769 696 1815 836
rect 1983 682 2029 728
rect 2187 699 2233 839
rect 2391 682 2437 728
rect 2595 683 2641 823
rect 2799 699 2845 839
rect 3003 699 3049 839
rect 3207 683 3253 823
rect 1185 589 1231 635
<< polysilicon >>
rect 608 944 2566 984
rect 134 852 234 896
rect 404 852 504 896
rect 608 852 708 944
rect 816 852 916 896
rect 1056 852 1156 896
rect 1436 852 1536 896
rect 1640 852 1740 896
rect 2058 852 2158 896
rect 2262 852 2362 896
rect 2466 852 2566 944
rect 2670 944 3178 984
rect 2670 852 2770 944
rect 2874 852 2974 896
rect 3078 852 3178 944
rect 134 500 234 669
rect 404 601 504 669
rect 404 588 537 601
rect 404 542 478 588
rect 524 542 537 588
rect 404 529 537 542
rect 134 454 147 500
rect 193 454 234 500
rect 608 481 708 669
rect 134 332 234 454
rect 348 441 708 481
rect 816 500 916 669
rect 816 454 829 500
rect 875 454 916 500
rect 124 288 244 332
rect 348 288 468 441
rect 572 380 692 393
rect 572 334 585 380
rect 631 334 692 380
rect 572 288 692 334
rect 816 332 916 454
rect 1056 415 1156 576
rect 1436 521 1536 669
rect 1640 628 1740 669
rect 1640 582 1681 628
rect 1727 609 1740 628
rect 2058 625 2158 669
rect 2058 609 2138 625
rect 1727 582 2138 609
rect 1640 569 2138 582
rect 1436 481 1690 521
rect 1650 465 1690 481
rect 1650 452 1959 465
rect 1056 369 1069 415
rect 1115 380 1156 415
rect 1426 420 1594 433
rect 1115 369 1176 380
rect 1056 336 1176 369
rect 1426 374 1535 420
rect 1581 374 1594 420
rect 1426 361 1594 374
rect 1650 406 1900 452
rect 1946 406 1959 452
rect 1650 393 1959 406
rect 796 288 916 332
rect 1426 301 1546 361
rect 1650 301 1770 393
rect 2018 333 2138 569
rect 2262 500 2362 669
rect 2262 454 2275 500
rect 2321 454 2362 500
rect 2262 377 2362 454
rect 2466 513 2566 669
rect 2670 625 2770 669
rect 2874 625 2974 669
rect 3078 625 3178 669
rect 2934 513 2974 625
rect 2466 500 2886 513
rect 2466 454 2827 500
rect 2873 454 2886 500
rect 2466 441 2886 454
rect 2934 500 3034 513
rect 2934 454 2947 500
rect 2993 454 3034 500
rect 2242 333 2362 377
rect 2466 333 2586 377
rect 2690 333 2810 441
rect 2934 377 3034 454
rect 2914 333 3034 377
rect 3138 377 3178 625
rect 3138 333 3258 377
rect 124 112 244 156
rect 348 112 468 156
rect 572 112 692 156
rect 796 112 916 156
rect 1056 112 1176 156
rect 1426 125 1546 169
rect 1650 125 1770 169
rect 2018 157 2138 201
rect 2242 157 2362 201
rect 652 64 692 112
rect 2466 64 2586 201
rect 2690 157 2810 201
rect 2914 157 3034 201
rect 3138 157 3258 201
rect 3138 64 3178 157
rect 652 24 3178 64
<< polycontact >>
rect 478 542 524 588
rect 147 454 193 500
rect 829 454 875 500
rect 585 334 631 380
rect 1681 582 1727 628
rect 1069 369 1115 415
rect 1535 374 1581 420
rect 1900 406 1946 452
rect 2275 454 2321 500
rect 2827 454 2873 500
rect 2947 454 2993 500
<< metal1 >>
rect 0 918 3472 1098
rect 59 839 105 918
rect 59 688 105 699
rect 273 823 319 834
rect 533 823 899 834
rect 142 500 194 542
rect 142 454 147 500
rect 193 454 194 500
rect 142 354 194 454
rect 49 275 95 286
rect 49 90 95 229
rect 273 275 319 683
rect 386 683 533 691
rect 579 788 899 823
rect 386 645 579 683
rect 721 728 783 739
rect 721 682 737 728
rect 721 671 783 682
rect 853 727 899 788
rect 945 830 991 918
rect 1769 836 2141 847
rect 945 773 991 784
rect 1361 823 1407 834
rect 853 683 1361 727
rect 853 681 1407 683
rect 1351 672 1407 681
rect 1565 823 1611 834
rect 1815 801 2141 836
rect 1815 696 1854 801
rect 1769 685 1854 696
rect 386 275 432 645
rect 478 588 530 599
rect 524 542 530 588
rect 478 380 530 542
rect 478 334 585 380
rect 631 334 642 380
rect 721 275 767 671
rect 1150 589 1185 635
rect 1231 589 1251 635
rect 814 500 875 542
rect 814 454 829 500
rect 1150 466 1251 589
rect 814 354 875 454
rect 1058 415 1115 426
rect 1058 369 1069 415
rect 1058 358 1115 369
rect 386 229 497 275
rect 543 229 554 275
rect 273 218 319 229
rect 721 218 767 229
rect 945 275 991 286
rect 945 90 991 229
rect 1058 185 1104 358
rect 1205 318 1251 466
rect 1150 299 1251 318
rect 1150 253 1205 299
rect 1150 242 1251 253
rect 1351 288 1397 672
rect 1565 523 1611 683
rect 1351 231 1397 242
rect 1443 477 1611 523
rect 1681 628 1762 639
rect 1727 582 1762 628
rect 1443 185 1489 477
rect 1681 431 1762 582
rect 1535 420 1762 431
rect 1581 374 1762 420
rect 1535 354 1762 374
rect 1808 286 1854 685
rect 1983 728 2029 739
rect 1983 463 2029 682
rect 2095 642 2141 801
rect 2187 839 2233 918
rect 2799 839 2845 850
rect 2187 688 2233 699
rect 2279 823 2661 834
rect 2279 788 2595 823
rect 2279 642 2325 788
rect 2095 596 2325 642
rect 2391 728 2437 739
rect 1799 275 1854 286
rect 1575 258 1621 269
rect 1845 229 1854 275
rect 1799 218 1854 229
rect 1900 452 2029 463
rect 1946 406 2029 452
rect 1900 275 2029 406
rect 2270 500 2322 542
rect 2270 454 2275 500
rect 2321 454 2322 500
rect 2270 354 2322 454
rect 1900 229 1943 275
rect 1989 229 2029 275
rect 1900 218 2029 229
rect 2167 275 2213 286
rect 1575 185 1621 212
rect 1058 139 1621 185
rect 2167 90 2213 229
rect 2391 275 2437 682
rect 2391 218 2437 229
rect 2641 683 2661 823
rect 2799 695 2845 699
rect 2595 275 2661 683
rect 2595 229 2615 275
rect 2735 649 2845 695
rect 3003 839 3049 918
rect 3003 688 3049 699
rect 3207 823 3253 834
rect 2735 275 2781 649
rect 3207 603 3253 683
rect 2827 557 3333 603
rect 2827 500 2873 557
rect 2827 443 2873 454
rect 2942 500 2994 511
rect 2942 454 2947 500
rect 2993 454 2994 500
rect 2735 229 2839 275
rect 2885 229 2896 275
rect 2942 242 2994 454
rect 3063 275 3109 286
rect 2595 218 2661 229
rect 3063 90 3109 229
rect 3287 275 3333 557
rect 3287 218 3333 229
rect 0 -90 3472 90
<< labels >>
flabel metal1 s 2942 242 2994 511 0 FreeSans 200 0 0 0 I0
port 1 nsew default input
flabel metal1 s 2270 354 2322 542 0 FreeSans 200 0 0 0 I1
port 2 nsew default input
flabel metal1 s 142 354 194 542 0 FreeSans 200 0 0 0 I2
port 3 nsew default input
flabel metal1 s 814 354 875 542 0 FreeSans 200 0 0 0 I3
port 4 nsew default input
flabel metal1 s 478 380 530 599 0 FreeSans 200 0 0 0 S0
port 5 nsew default input
flabel metal1 s 1681 431 1762 639 0 FreeSans 200 0 0 0 S1
port 6 nsew default input
flabel metal1 s 0 918 3472 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 3063 90 3109 286 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1150 466 1251 635 0 FreeSans 200 0 0 0 Z
port 7 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 478 334 642 380 1 S0
port 5 nsew default input
rlabel metal1 s 1535 354 1762 431 1 S1
port 6 nsew default input
rlabel metal1 s 1205 318 1251 466 1 Z
port 7 nsew default output
rlabel metal1 s 1150 242 1251 318 1 Z
port 7 nsew default output
rlabel metal1 s 3003 773 3049 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2187 773 2233 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 945 773 991 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 59 773 105 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3003 688 3049 773 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2187 688 2233 773 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 59 688 105 773 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2167 90 2213 286 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 945 90 991 286 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 49 90 95 286 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3472 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 1008
string GDS_END 14256
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 5716
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
