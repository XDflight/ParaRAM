magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal3 >>
rect 0 69639 200 69678
rect 800 69639 1000 69678
rect 0 69629 1000 69639
rect 0 69573 94 69629
rect 150 69573 218 69629
rect 274 69573 342 69629
rect 398 69573 466 69629
rect 522 69573 590 69629
rect 646 69573 714 69629
rect 770 69573 838 69629
rect 894 69573 1000 69629
rect 0 69505 1000 69573
rect 0 69449 94 69505
rect 150 69449 218 69505
rect 274 69449 342 69505
rect 398 69449 466 69505
rect 522 69449 590 69505
rect 646 69449 714 69505
rect 770 69449 838 69505
rect 894 69449 1000 69505
rect 0 69381 1000 69449
rect 0 69325 94 69381
rect 150 69325 218 69381
rect 274 69325 342 69381
rect 398 69325 466 69381
rect 522 69325 590 69381
rect 646 69325 714 69381
rect 770 69325 838 69381
rect 894 69325 1000 69381
rect 0 69257 1000 69325
rect 0 69201 94 69257
rect 150 69201 218 69257
rect 274 69201 342 69257
rect 398 69201 466 69257
rect 522 69201 590 69257
rect 646 69201 714 69257
rect 770 69201 838 69257
rect 894 69201 1000 69257
rect 0 69133 1000 69201
rect 0 69077 94 69133
rect 150 69077 218 69133
rect 274 69077 342 69133
rect 398 69077 466 69133
rect 522 69077 590 69133
rect 646 69077 714 69133
rect 770 69077 838 69133
rect 894 69077 1000 69133
rect 0 69009 1000 69077
rect 0 68953 94 69009
rect 150 68953 218 69009
rect 274 68953 342 69009
rect 398 68953 466 69009
rect 522 68953 590 69009
rect 646 68953 714 69009
rect 770 68953 838 69009
rect 894 68953 1000 69009
rect 0 68885 1000 68953
rect 0 68829 94 68885
rect 150 68829 218 68885
rect 274 68829 342 68885
rect 398 68829 466 68885
rect 522 68829 590 68885
rect 646 68829 714 68885
rect 770 68829 838 68885
rect 894 68829 1000 68885
rect 0 68761 1000 68829
rect 0 68705 94 68761
rect 150 68705 218 68761
rect 274 68705 342 68761
rect 398 68705 466 68761
rect 522 68705 590 68761
rect 646 68705 714 68761
rect 770 68705 838 68761
rect 894 68705 1000 68761
rect 0 68637 1000 68705
rect 0 68581 94 68637
rect 150 68581 218 68637
rect 274 68581 342 68637
rect 398 68581 466 68637
rect 522 68581 590 68637
rect 646 68581 714 68637
rect 770 68581 838 68637
rect 894 68581 1000 68637
rect 0 68513 1000 68581
rect 0 68457 94 68513
rect 150 68457 218 68513
rect 274 68457 342 68513
rect 398 68457 466 68513
rect 522 68457 590 68513
rect 646 68457 714 68513
rect 770 68457 838 68513
rect 894 68457 1000 68513
rect 0 68447 1000 68457
rect 0 68400 200 68447
rect 800 68400 1000 68447
rect 0 68094 200 68200
rect 800 68094 1000 68200
rect 0 68084 1000 68094
rect 0 68028 94 68084
rect 150 68028 218 68084
rect 274 68028 342 68084
rect 398 68028 466 68084
rect 522 68028 590 68084
rect 646 68028 714 68084
rect 770 68028 838 68084
rect 894 68028 1000 68084
rect 0 67960 1000 68028
rect 0 67904 94 67960
rect 150 67904 218 67960
rect 274 67904 342 67960
rect 398 67904 466 67960
rect 522 67904 590 67960
rect 646 67904 714 67960
rect 770 67904 838 67960
rect 894 67904 1000 67960
rect 0 67836 1000 67904
rect 0 67780 94 67836
rect 150 67780 218 67836
rect 274 67780 342 67836
rect 398 67780 466 67836
rect 522 67780 590 67836
rect 646 67780 714 67836
rect 770 67780 838 67836
rect 894 67780 1000 67836
rect 0 67712 1000 67780
rect 0 67656 94 67712
rect 150 67656 218 67712
rect 274 67656 342 67712
rect 398 67656 466 67712
rect 522 67656 590 67712
rect 646 67656 714 67712
rect 770 67656 838 67712
rect 894 67656 1000 67712
rect 0 67588 1000 67656
rect 0 67532 94 67588
rect 150 67532 218 67588
rect 274 67532 342 67588
rect 398 67532 466 67588
rect 522 67532 590 67588
rect 646 67532 714 67588
rect 770 67532 838 67588
rect 894 67532 1000 67588
rect 0 67464 1000 67532
rect 0 67408 94 67464
rect 150 67408 218 67464
rect 274 67408 342 67464
rect 398 67408 466 67464
rect 522 67408 590 67464
rect 646 67408 714 67464
rect 770 67408 838 67464
rect 894 67408 1000 67464
rect 0 67340 1000 67408
rect 0 67284 94 67340
rect 150 67284 218 67340
rect 274 67284 342 67340
rect 398 67284 466 67340
rect 522 67284 590 67340
rect 646 67284 714 67340
rect 770 67284 838 67340
rect 894 67284 1000 67340
rect 0 67216 1000 67284
rect 0 67160 94 67216
rect 150 67160 218 67216
rect 274 67160 342 67216
rect 398 67160 466 67216
rect 522 67160 590 67216
rect 646 67160 714 67216
rect 770 67160 838 67216
rect 894 67160 1000 67216
rect 0 67092 1000 67160
rect 0 67036 94 67092
rect 150 67036 218 67092
rect 274 67036 342 67092
rect 398 67036 466 67092
rect 522 67036 590 67092
rect 646 67036 714 67092
rect 770 67036 838 67092
rect 894 67036 1000 67092
rect 0 66968 1000 67036
rect 0 66912 94 66968
rect 150 66912 218 66968
rect 274 66912 342 66968
rect 398 66912 466 66968
rect 522 66912 590 66968
rect 646 66912 714 66968
rect 770 66912 838 66968
rect 894 66912 1000 66968
rect 0 66902 1000 66912
rect 0 66800 200 66902
rect 800 66800 1000 66902
rect 0 66487 200 66600
rect 800 66487 1000 66600
rect 0 66477 1000 66487
rect 0 66421 94 66477
rect 150 66421 218 66477
rect 274 66421 342 66477
rect 398 66421 466 66477
rect 522 66421 590 66477
rect 646 66421 714 66477
rect 770 66421 838 66477
rect 894 66421 1000 66477
rect 0 66353 1000 66421
rect 0 66297 94 66353
rect 150 66297 218 66353
rect 274 66297 342 66353
rect 398 66297 466 66353
rect 522 66297 590 66353
rect 646 66297 714 66353
rect 770 66297 838 66353
rect 894 66297 1000 66353
rect 0 66229 1000 66297
rect 0 66173 94 66229
rect 150 66173 218 66229
rect 274 66173 342 66229
rect 398 66173 466 66229
rect 522 66173 590 66229
rect 646 66173 714 66229
rect 770 66173 838 66229
rect 894 66173 1000 66229
rect 0 66105 1000 66173
rect 0 66049 94 66105
rect 150 66049 218 66105
rect 274 66049 342 66105
rect 398 66049 466 66105
rect 522 66049 590 66105
rect 646 66049 714 66105
rect 770 66049 838 66105
rect 894 66049 1000 66105
rect 0 65981 1000 66049
rect 0 65925 94 65981
rect 150 65925 218 65981
rect 274 65925 342 65981
rect 398 65925 466 65981
rect 522 65925 590 65981
rect 646 65925 714 65981
rect 770 65925 838 65981
rect 894 65925 1000 65981
rect 0 65857 1000 65925
rect 0 65801 94 65857
rect 150 65801 218 65857
rect 274 65801 342 65857
rect 398 65801 466 65857
rect 522 65801 590 65857
rect 646 65801 714 65857
rect 770 65801 838 65857
rect 894 65801 1000 65857
rect 0 65733 1000 65801
rect 0 65677 94 65733
rect 150 65677 218 65733
rect 274 65677 342 65733
rect 398 65677 466 65733
rect 522 65677 590 65733
rect 646 65677 714 65733
rect 770 65677 838 65733
rect 894 65677 1000 65733
rect 0 65609 1000 65677
rect 0 65553 94 65609
rect 150 65553 218 65609
rect 274 65553 342 65609
rect 398 65553 466 65609
rect 522 65553 590 65609
rect 646 65553 714 65609
rect 770 65553 838 65609
rect 894 65553 1000 65609
rect 0 65485 1000 65553
rect 0 65429 94 65485
rect 150 65429 218 65485
rect 274 65429 342 65485
rect 398 65429 466 65485
rect 522 65429 590 65485
rect 646 65429 714 65485
rect 770 65429 838 65485
rect 894 65429 1000 65485
rect 0 65361 1000 65429
rect 0 65305 94 65361
rect 150 65305 218 65361
rect 274 65305 342 65361
rect 398 65305 466 65361
rect 522 65305 590 65361
rect 646 65305 714 65361
rect 770 65305 838 65361
rect 894 65305 1000 65361
rect 0 65295 1000 65305
rect 0 65200 200 65295
rect 800 65200 1000 65295
rect 0 64896 200 65000
rect 800 64896 1000 65000
rect 0 64886 1000 64896
rect 0 64830 94 64886
rect 150 64830 218 64886
rect 274 64830 342 64886
rect 398 64830 466 64886
rect 522 64830 590 64886
rect 646 64830 714 64886
rect 770 64830 838 64886
rect 894 64830 1000 64886
rect 0 64762 1000 64830
rect 0 64706 94 64762
rect 150 64706 218 64762
rect 274 64706 342 64762
rect 398 64706 466 64762
rect 522 64706 590 64762
rect 646 64706 714 64762
rect 770 64706 838 64762
rect 894 64706 1000 64762
rect 0 64638 1000 64706
rect 0 64582 94 64638
rect 150 64582 218 64638
rect 274 64582 342 64638
rect 398 64582 466 64638
rect 522 64582 590 64638
rect 646 64582 714 64638
rect 770 64582 838 64638
rect 894 64582 1000 64638
rect 0 64514 1000 64582
rect 0 64458 94 64514
rect 150 64458 218 64514
rect 274 64458 342 64514
rect 398 64458 466 64514
rect 522 64458 590 64514
rect 646 64458 714 64514
rect 770 64458 838 64514
rect 894 64458 1000 64514
rect 0 64390 1000 64458
rect 0 64334 94 64390
rect 150 64334 218 64390
rect 274 64334 342 64390
rect 398 64334 466 64390
rect 522 64334 590 64390
rect 646 64334 714 64390
rect 770 64334 838 64390
rect 894 64334 1000 64390
rect 0 64266 1000 64334
rect 0 64210 94 64266
rect 150 64210 218 64266
rect 274 64210 342 64266
rect 398 64210 466 64266
rect 522 64210 590 64266
rect 646 64210 714 64266
rect 770 64210 838 64266
rect 894 64210 1000 64266
rect 0 64142 1000 64210
rect 0 64086 94 64142
rect 150 64086 218 64142
rect 274 64086 342 64142
rect 398 64086 466 64142
rect 522 64086 590 64142
rect 646 64086 714 64142
rect 770 64086 838 64142
rect 894 64086 1000 64142
rect 0 64018 1000 64086
rect 0 63962 94 64018
rect 150 63962 218 64018
rect 274 63962 342 64018
rect 398 63962 466 64018
rect 522 63962 590 64018
rect 646 63962 714 64018
rect 770 63962 838 64018
rect 894 63962 1000 64018
rect 0 63894 1000 63962
rect 0 63838 94 63894
rect 150 63838 218 63894
rect 274 63838 342 63894
rect 398 63838 466 63894
rect 522 63838 590 63894
rect 646 63838 714 63894
rect 770 63838 838 63894
rect 894 63838 1000 63894
rect 0 63770 1000 63838
rect 0 63714 94 63770
rect 150 63714 218 63770
rect 274 63714 342 63770
rect 398 63714 466 63770
rect 522 63714 590 63770
rect 646 63714 714 63770
rect 770 63714 838 63770
rect 894 63714 1000 63770
rect 0 63704 1000 63714
rect 0 63600 200 63704
rect 800 63600 1000 63704
rect 0 63290 200 63400
rect 800 63290 1000 63400
rect 0 63280 1000 63290
rect 0 63224 94 63280
rect 150 63224 218 63280
rect 274 63224 342 63280
rect 398 63224 466 63280
rect 522 63224 590 63280
rect 646 63224 714 63280
rect 770 63224 838 63280
rect 894 63224 1000 63280
rect 0 63156 1000 63224
rect 0 63100 94 63156
rect 150 63100 218 63156
rect 274 63100 342 63156
rect 398 63100 466 63156
rect 522 63100 590 63156
rect 646 63100 714 63156
rect 770 63100 838 63156
rect 894 63100 1000 63156
rect 0 63032 1000 63100
rect 0 62976 94 63032
rect 150 62976 218 63032
rect 274 62976 342 63032
rect 398 62976 466 63032
rect 522 62976 590 63032
rect 646 62976 714 63032
rect 770 62976 838 63032
rect 894 62976 1000 63032
rect 0 62908 1000 62976
rect 0 62852 94 62908
rect 150 62852 218 62908
rect 274 62852 342 62908
rect 398 62852 466 62908
rect 522 62852 590 62908
rect 646 62852 714 62908
rect 770 62852 838 62908
rect 894 62852 1000 62908
rect 0 62784 1000 62852
rect 0 62728 94 62784
rect 150 62728 218 62784
rect 274 62728 342 62784
rect 398 62728 466 62784
rect 522 62728 590 62784
rect 646 62728 714 62784
rect 770 62728 838 62784
rect 894 62728 1000 62784
rect 0 62660 1000 62728
rect 0 62604 94 62660
rect 150 62604 218 62660
rect 274 62604 342 62660
rect 398 62604 466 62660
rect 522 62604 590 62660
rect 646 62604 714 62660
rect 770 62604 838 62660
rect 894 62604 1000 62660
rect 0 62536 1000 62604
rect 0 62480 94 62536
rect 150 62480 218 62536
rect 274 62480 342 62536
rect 398 62480 466 62536
rect 522 62480 590 62536
rect 646 62480 714 62536
rect 770 62480 838 62536
rect 894 62480 1000 62536
rect 0 62412 1000 62480
rect 0 62356 94 62412
rect 150 62356 218 62412
rect 274 62356 342 62412
rect 398 62356 466 62412
rect 522 62356 590 62412
rect 646 62356 714 62412
rect 770 62356 838 62412
rect 894 62356 1000 62412
rect 0 62288 1000 62356
rect 0 62232 94 62288
rect 150 62232 218 62288
rect 274 62232 342 62288
rect 398 62232 466 62288
rect 522 62232 590 62288
rect 646 62232 714 62288
rect 770 62232 838 62288
rect 894 62232 1000 62288
rect 0 62164 1000 62232
rect 0 62108 94 62164
rect 150 62108 218 62164
rect 274 62108 342 62164
rect 398 62108 466 62164
rect 522 62108 590 62164
rect 646 62108 714 62164
rect 770 62108 838 62164
rect 894 62108 1000 62164
rect 0 62098 1000 62108
rect 0 62000 200 62098
rect 800 62000 1000 62098
rect 0 61704 200 61800
rect 800 61704 1000 61800
rect 0 61694 1000 61704
rect 0 61638 94 61694
rect 150 61638 218 61694
rect 274 61638 342 61694
rect 398 61638 466 61694
rect 522 61638 590 61694
rect 646 61638 714 61694
rect 770 61638 838 61694
rect 894 61638 1000 61694
rect 0 61570 1000 61638
rect 0 61514 94 61570
rect 150 61514 218 61570
rect 274 61514 342 61570
rect 398 61514 466 61570
rect 522 61514 590 61570
rect 646 61514 714 61570
rect 770 61514 838 61570
rect 894 61514 1000 61570
rect 0 61446 1000 61514
rect 0 61390 94 61446
rect 150 61390 218 61446
rect 274 61390 342 61446
rect 398 61390 466 61446
rect 522 61390 590 61446
rect 646 61390 714 61446
rect 770 61390 838 61446
rect 894 61390 1000 61446
rect 0 61322 1000 61390
rect 0 61266 94 61322
rect 150 61266 218 61322
rect 274 61266 342 61322
rect 398 61266 466 61322
rect 522 61266 590 61322
rect 646 61266 714 61322
rect 770 61266 838 61322
rect 894 61266 1000 61322
rect 0 61198 1000 61266
rect 0 61142 94 61198
rect 150 61142 218 61198
rect 274 61142 342 61198
rect 398 61142 466 61198
rect 522 61142 590 61198
rect 646 61142 714 61198
rect 770 61142 838 61198
rect 894 61142 1000 61198
rect 0 61074 1000 61142
rect 0 61018 94 61074
rect 150 61018 218 61074
rect 274 61018 342 61074
rect 398 61018 466 61074
rect 522 61018 590 61074
rect 646 61018 714 61074
rect 770 61018 838 61074
rect 894 61018 1000 61074
rect 0 60950 1000 61018
rect 0 60894 94 60950
rect 150 60894 218 60950
rect 274 60894 342 60950
rect 398 60894 466 60950
rect 522 60894 590 60950
rect 646 60894 714 60950
rect 770 60894 838 60950
rect 894 60894 1000 60950
rect 0 60826 1000 60894
rect 0 60770 94 60826
rect 150 60770 218 60826
rect 274 60770 342 60826
rect 398 60770 466 60826
rect 522 60770 590 60826
rect 646 60770 714 60826
rect 770 60770 838 60826
rect 894 60770 1000 60826
rect 0 60702 1000 60770
rect 0 60646 94 60702
rect 150 60646 218 60702
rect 274 60646 342 60702
rect 398 60646 466 60702
rect 522 60646 590 60702
rect 646 60646 714 60702
rect 770 60646 838 60702
rect 894 60646 1000 60702
rect 0 60578 1000 60646
rect 0 60522 94 60578
rect 150 60522 218 60578
rect 274 60522 342 60578
rect 398 60522 466 60578
rect 522 60522 590 60578
rect 646 60522 714 60578
rect 770 60522 838 60578
rect 894 60522 1000 60578
rect 0 60512 1000 60522
rect 0 60400 200 60512
rect 800 60400 1000 60512
rect 0 60112 200 60200
rect 800 60112 1000 60200
rect 0 60102 1000 60112
rect 0 60046 94 60102
rect 150 60046 218 60102
rect 274 60046 342 60102
rect 398 60046 466 60102
rect 522 60046 590 60102
rect 646 60046 714 60102
rect 770 60046 838 60102
rect 894 60046 1000 60102
rect 0 59978 1000 60046
rect 0 59922 94 59978
rect 150 59922 218 59978
rect 274 59922 342 59978
rect 398 59922 466 59978
rect 522 59922 590 59978
rect 646 59922 714 59978
rect 770 59922 838 59978
rect 894 59922 1000 59978
rect 0 59854 1000 59922
rect 0 59798 94 59854
rect 150 59798 218 59854
rect 274 59798 342 59854
rect 398 59798 466 59854
rect 522 59798 590 59854
rect 646 59798 714 59854
rect 770 59798 838 59854
rect 894 59798 1000 59854
rect 0 59730 1000 59798
rect 0 59674 94 59730
rect 150 59674 218 59730
rect 274 59674 342 59730
rect 398 59674 466 59730
rect 522 59674 590 59730
rect 646 59674 714 59730
rect 770 59674 838 59730
rect 894 59674 1000 59730
rect 0 59606 1000 59674
rect 0 59550 94 59606
rect 150 59550 218 59606
rect 274 59550 342 59606
rect 398 59550 466 59606
rect 522 59550 590 59606
rect 646 59550 714 59606
rect 770 59550 838 59606
rect 894 59550 1000 59606
rect 0 59482 1000 59550
rect 0 59426 94 59482
rect 150 59426 218 59482
rect 274 59426 342 59482
rect 398 59426 466 59482
rect 522 59426 590 59482
rect 646 59426 714 59482
rect 770 59426 838 59482
rect 894 59426 1000 59482
rect 0 59358 1000 59426
rect 0 59302 94 59358
rect 150 59302 218 59358
rect 274 59302 342 59358
rect 398 59302 466 59358
rect 522 59302 590 59358
rect 646 59302 714 59358
rect 770 59302 838 59358
rect 894 59302 1000 59358
rect 0 59234 1000 59302
rect 0 59178 94 59234
rect 150 59178 218 59234
rect 274 59178 342 59234
rect 398 59178 466 59234
rect 522 59178 590 59234
rect 646 59178 714 59234
rect 770 59178 838 59234
rect 894 59178 1000 59234
rect 0 59110 1000 59178
rect 0 59054 94 59110
rect 150 59054 218 59110
rect 274 59054 342 59110
rect 398 59054 466 59110
rect 522 59054 590 59110
rect 646 59054 714 59110
rect 770 59054 838 59110
rect 894 59054 1000 59110
rect 0 58986 1000 59054
rect 0 58930 94 58986
rect 150 58930 218 58986
rect 274 58930 342 58986
rect 398 58930 466 58986
rect 522 58930 590 58986
rect 646 58930 714 58986
rect 770 58930 838 58986
rect 894 58930 1000 58986
rect 0 58920 1000 58930
rect 0 58800 200 58920
rect 800 58800 1000 58920
rect 0 58495 200 58600
rect 800 58495 1000 58600
rect 0 58485 1000 58495
rect 0 58429 94 58485
rect 150 58429 218 58485
rect 274 58429 342 58485
rect 398 58429 466 58485
rect 522 58429 590 58485
rect 646 58429 714 58485
rect 770 58429 838 58485
rect 894 58429 1000 58485
rect 0 58361 1000 58429
rect 0 58305 94 58361
rect 150 58305 218 58361
rect 274 58305 342 58361
rect 398 58305 466 58361
rect 522 58305 590 58361
rect 646 58305 714 58361
rect 770 58305 838 58361
rect 894 58305 1000 58361
rect 0 58237 1000 58305
rect 0 58181 94 58237
rect 150 58181 218 58237
rect 274 58181 342 58237
rect 398 58181 466 58237
rect 522 58181 590 58237
rect 646 58181 714 58237
rect 770 58181 838 58237
rect 894 58181 1000 58237
rect 0 58113 1000 58181
rect 0 58057 94 58113
rect 150 58057 218 58113
rect 274 58057 342 58113
rect 398 58057 466 58113
rect 522 58057 590 58113
rect 646 58057 714 58113
rect 770 58057 838 58113
rect 894 58057 1000 58113
rect 0 57989 1000 58057
rect 0 57933 94 57989
rect 150 57933 218 57989
rect 274 57933 342 57989
rect 398 57933 466 57989
rect 522 57933 590 57989
rect 646 57933 714 57989
rect 770 57933 838 57989
rect 894 57933 1000 57989
rect 0 57865 1000 57933
rect 0 57809 94 57865
rect 150 57809 218 57865
rect 274 57809 342 57865
rect 398 57809 466 57865
rect 522 57809 590 57865
rect 646 57809 714 57865
rect 770 57809 838 57865
rect 894 57809 1000 57865
rect 0 57741 1000 57809
rect 0 57685 94 57741
rect 150 57685 218 57741
rect 274 57685 342 57741
rect 398 57685 466 57741
rect 522 57685 590 57741
rect 646 57685 714 57741
rect 770 57685 838 57741
rect 894 57685 1000 57741
rect 0 57617 1000 57685
rect 0 57561 94 57617
rect 150 57561 218 57617
rect 274 57561 342 57617
rect 398 57561 466 57617
rect 522 57561 590 57617
rect 646 57561 714 57617
rect 770 57561 838 57617
rect 894 57561 1000 57617
rect 0 57493 1000 57561
rect 0 57437 94 57493
rect 150 57437 218 57493
rect 274 57437 342 57493
rect 398 57437 466 57493
rect 522 57437 590 57493
rect 646 57437 714 57493
rect 770 57437 838 57493
rect 894 57437 1000 57493
rect 0 57369 1000 57437
rect 0 57313 94 57369
rect 150 57313 218 57369
rect 274 57313 342 57369
rect 398 57313 466 57369
rect 522 57313 590 57369
rect 646 57313 714 57369
rect 770 57313 838 57369
rect 894 57313 1000 57369
rect 0 57303 1000 57313
rect 0 57200 200 57303
rect 800 57200 1000 57303
rect 0 56902 200 57000
rect 800 56902 1000 57000
rect 0 56892 1000 56902
rect 0 56836 94 56892
rect 150 56836 218 56892
rect 274 56836 342 56892
rect 398 56836 466 56892
rect 522 56836 590 56892
rect 646 56836 714 56892
rect 770 56836 838 56892
rect 894 56836 1000 56892
rect 0 56768 1000 56836
rect 0 56712 94 56768
rect 150 56712 218 56768
rect 274 56712 342 56768
rect 398 56712 466 56768
rect 522 56712 590 56768
rect 646 56712 714 56768
rect 770 56712 838 56768
rect 894 56712 1000 56768
rect 0 56644 1000 56712
rect 0 56588 94 56644
rect 150 56588 218 56644
rect 274 56588 342 56644
rect 398 56588 466 56644
rect 522 56588 590 56644
rect 646 56588 714 56644
rect 770 56588 838 56644
rect 894 56588 1000 56644
rect 0 56520 1000 56588
rect 0 56464 94 56520
rect 150 56464 218 56520
rect 274 56464 342 56520
rect 398 56464 466 56520
rect 522 56464 590 56520
rect 646 56464 714 56520
rect 770 56464 838 56520
rect 894 56464 1000 56520
rect 0 56396 1000 56464
rect 0 56340 94 56396
rect 150 56340 218 56396
rect 274 56340 342 56396
rect 398 56340 466 56396
rect 522 56340 590 56396
rect 646 56340 714 56396
rect 770 56340 838 56396
rect 894 56340 1000 56396
rect 0 56272 1000 56340
rect 0 56216 94 56272
rect 150 56216 218 56272
rect 274 56216 342 56272
rect 398 56216 466 56272
rect 522 56216 590 56272
rect 646 56216 714 56272
rect 770 56216 838 56272
rect 894 56216 1000 56272
rect 0 56148 1000 56216
rect 0 56092 94 56148
rect 150 56092 218 56148
rect 274 56092 342 56148
rect 398 56092 466 56148
rect 522 56092 590 56148
rect 646 56092 714 56148
rect 770 56092 838 56148
rect 894 56092 1000 56148
rect 0 56024 1000 56092
rect 0 55968 94 56024
rect 150 55968 218 56024
rect 274 55968 342 56024
rect 398 55968 466 56024
rect 522 55968 590 56024
rect 646 55968 714 56024
rect 770 55968 838 56024
rect 894 55968 1000 56024
rect 0 55900 1000 55968
rect 0 55844 94 55900
rect 150 55844 218 55900
rect 274 55844 342 55900
rect 398 55844 466 55900
rect 522 55844 590 55900
rect 646 55844 714 55900
rect 770 55844 838 55900
rect 894 55844 1000 55900
rect 0 55776 1000 55844
rect 0 55720 94 55776
rect 150 55720 218 55776
rect 274 55720 342 55776
rect 398 55720 466 55776
rect 522 55720 590 55776
rect 646 55720 714 55776
rect 770 55720 838 55776
rect 894 55720 1000 55776
rect 0 55710 1000 55720
rect 0 55600 200 55710
rect 800 55600 1000 55710
rect 0 55298 200 55400
rect 800 55298 1000 55400
rect 0 55288 1000 55298
rect 0 55232 94 55288
rect 150 55232 218 55288
rect 274 55232 342 55288
rect 398 55232 466 55288
rect 522 55232 590 55288
rect 646 55232 714 55288
rect 770 55232 838 55288
rect 894 55232 1000 55288
rect 0 55164 1000 55232
rect 0 55108 94 55164
rect 150 55108 218 55164
rect 274 55108 342 55164
rect 398 55108 466 55164
rect 522 55108 590 55164
rect 646 55108 714 55164
rect 770 55108 838 55164
rect 894 55108 1000 55164
rect 0 55040 1000 55108
rect 0 54984 94 55040
rect 150 54984 218 55040
rect 274 54984 342 55040
rect 398 54984 466 55040
rect 522 54984 590 55040
rect 646 54984 714 55040
rect 770 54984 838 55040
rect 894 54984 1000 55040
rect 0 54916 1000 54984
rect 0 54860 94 54916
rect 150 54860 218 54916
rect 274 54860 342 54916
rect 398 54860 466 54916
rect 522 54860 590 54916
rect 646 54860 714 54916
rect 770 54860 838 54916
rect 894 54860 1000 54916
rect 0 54792 1000 54860
rect 0 54736 94 54792
rect 150 54736 218 54792
rect 274 54736 342 54792
rect 398 54736 466 54792
rect 522 54736 590 54792
rect 646 54736 714 54792
rect 770 54736 838 54792
rect 894 54736 1000 54792
rect 0 54668 1000 54736
rect 0 54612 94 54668
rect 150 54612 218 54668
rect 274 54612 342 54668
rect 398 54612 466 54668
rect 522 54612 590 54668
rect 646 54612 714 54668
rect 770 54612 838 54668
rect 894 54612 1000 54668
rect 0 54544 1000 54612
rect 0 54488 94 54544
rect 150 54488 218 54544
rect 274 54488 342 54544
rect 398 54488 466 54544
rect 522 54488 590 54544
rect 646 54488 714 54544
rect 770 54488 838 54544
rect 894 54488 1000 54544
rect 0 54420 1000 54488
rect 0 54364 94 54420
rect 150 54364 218 54420
rect 274 54364 342 54420
rect 398 54364 466 54420
rect 522 54364 590 54420
rect 646 54364 714 54420
rect 770 54364 838 54420
rect 894 54364 1000 54420
rect 0 54296 1000 54364
rect 0 54240 94 54296
rect 150 54240 218 54296
rect 274 54240 342 54296
rect 398 54240 466 54296
rect 522 54240 590 54296
rect 646 54240 714 54296
rect 770 54240 838 54296
rect 894 54240 1000 54296
rect 0 54172 1000 54240
rect 0 54116 94 54172
rect 150 54116 218 54172
rect 274 54116 342 54172
rect 398 54116 466 54172
rect 522 54116 590 54172
rect 646 54116 714 54172
rect 770 54116 838 54172
rect 894 54116 1000 54172
rect 0 54106 1000 54116
rect 0 54000 200 54106
rect 800 54000 1000 54106
rect 0 53692 200 53800
rect 800 53692 1000 53800
rect 0 53682 1000 53692
rect 0 53626 94 53682
rect 150 53626 218 53682
rect 274 53626 342 53682
rect 398 53626 466 53682
rect 522 53626 590 53682
rect 646 53626 714 53682
rect 770 53626 838 53682
rect 894 53626 1000 53682
rect 0 53558 1000 53626
rect 0 53502 94 53558
rect 150 53502 218 53558
rect 274 53502 342 53558
rect 398 53502 466 53558
rect 522 53502 590 53558
rect 646 53502 714 53558
rect 770 53502 838 53558
rect 894 53502 1000 53558
rect 0 53434 1000 53502
rect 0 53378 94 53434
rect 150 53378 218 53434
rect 274 53378 342 53434
rect 398 53378 466 53434
rect 522 53378 590 53434
rect 646 53378 714 53434
rect 770 53378 838 53434
rect 894 53378 1000 53434
rect 0 53310 1000 53378
rect 0 53254 94 53310
rect 150 53254 218 53310
rect 274 53254 342 53310
rect 398 53254 466 53310
rect 522 53254 590 53310
rect 646 53254 714 53310
rect 770 53254 838 53310
rect 894 53254 1000 53310
rect 0 53186 1000 53254
rect 0 53130 94 53186
rect 150 53130 218 53186
rect 274 53130 342 53186
rect 398 53130 466 53186
rect 522 53130 590 53186
rect 646 53130 714 53186
rect 770 53130 838 53186
rect 894 53130 1000 53186
rect 0 53062 1000 53130
rect 0 53006 94 53062
rect 150 53006 218 53062
rect 274 53006 342 53062
rect 398 53006 466 53062
rect 522 53006 590 53062
rect 646 53006 714 53062
rect 770 53006 838 53062
rect 894 53006 1000 53062
rect 0 52938 1000 53006
rect 0 52882 94 52938
rect 150 52882 218 52938
rect 274 52882 342 52938
rect 398 52882 466 52938
rect 522 52882 590 52938
rect 646 52882 714 52938
rect 770 52882 838 52938
rect 894 52882 1000 52938
rect 0 52814 1000 52882
rect 0 52758 94 52814
rect 150 52758 218 52814
rect 274 52758 342 52814
rect 398 52758 466 52814
rect 522 52758 590 52814
rect 646 52758 714 52814
rect 770 52758 838 52814
rect 894 52758 1000 52814
rect 0 52690 1000 52758
rect 0 52634 94 52690
rect 150 52634 218 52690
rect 274 52634 342 52690
rect 398 52634 466 52690
rect 522 52634 590 52690
rect 646 52634 714 52690
rect 770 52634 838 52690
rect 894 52634 1000 52690
rect 0 52566 1000 52634
rect 0 52510 94 52566
rect 150 52510 218 52566
rect 274 52510 342 52566
rect 398 52510 466 52566
rect 522 52510 590 52566
rect 646 52510 714 52566
rect 770 52510 838 52566
rect 894 52510 1000 52566
rect 0 52500 1000 52510
rect 0 52400 200 52500
rect 800 52400 1000 52500
rect 0 52089 200 52200
rect 800 52089 1000 52200
rect 0 52079 1000 52089
rect 0 52023 94 52079
rect 150 52023 218 52079
rect 274 52023 342 52079
rect 398 52023 466 52079
rect 522 52023 590 52079
rect 646 52023 714 52079
rect 770 52023 838 52079
rect 894 52023 1000 52079
rect 0 51955 1000 52023
rect 0 51899 94 51955
rect 150 51899 218 51955
rect 274 51899 342 51955
rect 398 51899 466 51955
rect 522 51899 590 51955
rect 646 51899 714 51955
rect 770 51899 838 51955
rect 894 51899 1000 51955
rect 0 51831 1000 51899
rect 0 51775 94 51831
rect 150 51775 218 51831
rect 274 51775 342 51831
rect 398 51775 466 51831
rect 522 51775 590 51831
rect 646 51775 714 51831
rect 770 51775 838 51831
rect 894 51775 1000 51831
rect 0 51707 1000 51775
rect 0 51651 94 51707
rect 150 51651 218 51707
rect 274 51651 342 51707
rect 398 51651 466 51707
rect 522 51651 590 51707
rect 646 51651 714 51707
rect 770 51651 838 51707
rect 894 51651 1000 51707
rect 0 51583 1000 51651
rect 0 51527 94 51583
rect 150 51527 218 51583
rect 274 51527 342 51583
rect 398 51527 466 51583
rect 522 51527 590 51583
rect 646 51527 714 51583
rect 770 51527 838 51583
rect 894 51527 1000 51583
rect 0 51459 1000 51527
rect 0 51403 94 51459
rect 150 51403 218 51459
rect 274 51403 342 51459
rect 398 51403 466 51459
rect 522 51403 590 51459
rect 646 51403 714 51459
rect 770 51403 838 51459
rect 894 51403 1000 51459
rect 0 51335 1000 51403
rect 0 51279 94 51335
rect 150 51279 218 51335
rect 274 51279 342 51335
rect 398 51279 466 51335
rect 522 51279 590 51335
rect 646 51279 714 51335
rect 770 51279 838 51335
rect 894 51279 1000 51335
rect 0 51211 1000 51279
rect 0 51155 94 51211
rect 150 51155 218 51211
rect 274 51155 342 51211
rect 398 51155 466 51211
rect 522 51155 590 51211
rect 646 51155 714 51211
rect 770 51155 838 51211
rect 894 51155 1000 51211
rect 0 51087 1000 51155
rect 0 51031 94 51087
rect 150 51031 218 51087
rect 274 51031 342 51087
rect 398 51031 466 51087
rect 522 51031 590 51087
rect 646 51031 714 51087
rect 770 51031 838 51087
rect 894 51031 1000 51087
rect 0 50963 1000 51031
rect 0 50907 94 50963
rect 150 50907 218 50963
rect 274 50907 342 50963
rect 398 50907 466 50963
rect 522 50907 590 50963
rect 646 50907 714 50963
rect 770 50907 838 50963
rect 894 50907 1000 50963
rect 0 50897 1000 50907
rect 0 50800 200 50897
rect 800 50800 1000 50897
rect 0 50490 200 50600
rect 800 50490 1000 50600
rect 0 50480 1000 50490
rect 0 50424 95 50480
rect 151 50424 219 50480
rect 275 50424 343 50480
rect 399 50424 467 50480
rect 523 50424 591 50480
rect 647 50424 715 50480
rect 771 50424 839 50480
rect 895 50424 1000 50480
rect 0 50356 1000 50424
rect 0 50300 95 50356
rect 151 50300 219 50356
rect 275 50300 343 50356
rect 399 50300 467 50356
rect 523 50300 591 50356
rect 647 50300 715 50356
rect 771 50300 839 50356
rect 895 50300 1000 50356
rect 0 50232 1000 50300
rect 0 50176 95 50232
rect 151 50176 219 50232
rect 275 50176 343 50232
rect 399 50176 467 50232
rect 523 50176 591 50232
rect 647 50176 715 50232
rect 771 50176 839 50232
rect 895 50176 1000 50232
rect 0 50108 1000 50176
rect 0 50052 95 50108
rect 151 50052 219 50108
rect 275 50052 343 50108
rect 399 50052 467 50108
rect 523 50052 591 50108
rect 647 50052 715 50108
rect 771 50052 839 50108
rect 895 50052 1000 50108
rect 0 49984 1000 50052
rect 0 49928 95 49984
rect 151 49928 219 49984
rect 275 49928 343 49984
rect 399 49928 467 49984
rect 523 49928 591 49984
rect 647 49928 715 49984
rect 771 49928 839 49984
rect 895 49928 1000 49984
rect 0 49860 1000 49928
rect 0 49804 95 49860
rect 151 49804 219 49860
rect 275 49804 343 49860
rect 399 49804 467 49860
rect 523 49804 591 49860
rect 647 49804 715 49860
rect 771 49804 839 49860
rect 895 49804 1000 49860
rect 0 49736 1000 49804
rect 0 49680 95 49736
rect 151 49680 219 49736
rect 275 49680 343 49736
rect 399 49680 467 49736
rect 523 49680 591 49736
rect 647 49680 715 49736
rect 771 49680 839 49736
rect 895 49680 1000 49736
rect 0 49612 1000 49680
rect 0 49556 95 49612
rect 151 49556 219 49612
rect 275 49556 343 49612
rect 399 49556 467 49612
rect 523 49556 591 49612
rect 647 49556 715 49612
rect 771 49556 839 49612
rect 895 49556 1000 49612
rect 0 49488 1000 49556
rect 0 49432 95 49488
rect 151 49432 219 49488
rect 275 49432 343 49488
rect 399 49432 467 49488
rect 523 49432 591 49488
rect 647 49432 715 49488
rect 771 49432 839 49488
rect 895 49432 1000 49488
rect 0 49364 1000 49432
rect 0 49308 95 49364
rect 151 49308 219 49364
rect 275 49308 343 49364
rect 399 49308 467 49364
rect 523 49308 591 49364
rect 647 49308 715 49364
rect 771 49308 839 49364
rect 895 49308 1000 49364
rect 0 49298 1000 49308
rect 0 49200 200 49298
rect 800 49200 1000 49298
rect 0 48903 200 49000
rect 800 48903 1000 49000
rect 0 48893 1000 48903
rect 0 48837 94 48893
rect 150 48837 218 48893
rect 274 48837 342 48893
rect 398 48837 466 48893
rect 522 48837 590 48893
rect 646 48837 714 48893
rect 770 48837 838 48893
rect 894 48837 1000 48893
rect 0 48769 1000 48837
rect 0 48713 94 48769
rect 150 48713 218 48769
rect 274 48713 342 48769
rect 398 48713 466 48769
rect 522 48713 590 48769
rect 646 48713 714 48769
rect 770 48713 838 48769
rect 894 48713 1000 48769
rect 0 48645 1000 48713
rect 0 48589 94 48645
rect 150 48589 218 48645
rect 274 48589 342 48645
rect 398 48589 466 48645
rect 522 48589 590 48645
rect 646 48589 714 48645
rect 770 48589 838 48645
rect 894 48589 1000 48645
rect 0 48521 1000 48589
rect 0 48465 94 48521
rect 150 48465 218 48521
rect 274 48465 342 48521
rect 398 48465 466 48521
rect 522 48465 590 48521
rect 646 48465 714 48521
rect 770 48465 838 48521
rect 894 48465 1000 48521
rect 0 48397 1000 48465
rect 0 48341 94 48397
rect 150 48341 218 48397
rect 274 48341 342 48397
rect 398 48341 466 48397
rect 522 48341 590 48397
rect 646 48341 714 48397
rect 770 48341 838 48397
rect 894 48341 1000 48397
rect 0 48273 1000 48341
rect 0 48217 94 48273
rect 150 48217 218 48273
rect 274 48217 342 48273
rect 398 48217 466 48273
rect 522 48217 590 48273
rect 646 48217 714 48273
rect 770 48217 838 48273
rect 894 48217 1000 48273
rect 0 48149 1000 48217
rect 0 48093 94 48149
rect 150 48093 218 48149
rect 274 48093 342 48149
rect 398 48093 466 48149
rect 522 48093 590 48149
rect 646 48093 714 48149
rect 770 48093 838 48149
rect 894 48093 1000 48149
rect 0 48025 1000 48093
rect 0 47969 94 48025
rect 150 47969 218 48025
rect 274 47969 342 48025
rect 398 47969 466 48025
rect 522 47969 590 48025
rect 646 47969 714 48025
rect 770 47969 838 48025
rect 894 47969 1000 48025
rect 0 47901 1000 47969
rect 0 47845 94 47901
rect 150 47845 218 47901
rect 274 47845 342 47901
rect 398 47845 466 47901
rect 522 47845 590 47901
rect 646 47845 714 47901
rect 770 47845 838 47901
rect 894 47845 1000 47901
rect 0 47777 1000 47845
rect 0 47721 94 47777
rect 150 47721 218 47777
rect 274 47721 342 47777
rect 398 47721 466 47777
rect 522 47721 590 47777
rect 646 47721 714 47777
rect 770 47721 838 47777
rect 894 47721 1000 47777
rect 0 47653 1000 47721
rect 0 47597 94 47653
rect 150 47597 218 47653
rect 274 47597 342 47653
rect 398 47597 466 47653
rect 522 47597 590 47653
rect 646 47597 714 47653
rect 770 47597 838 47653
rect 894 47597 1000 47653
rect 0 47529 1000 47597
rect 0 47473 94 47529
rect 150 47473 218 47529
rect 274 47473 342 47529
rect 398 47473 466 47529
rect 522 47473 590 47529
rect 646 47473 714 47529
rect 770 47473 838 47529
rect 894 47473 1000 47529
rect 0 47405 1000 47473
rect 0 47349 94 47405
rect 150 47349 218 47405
rect 274 47349 342 47405
rect 398 47349 466 47405
rect 522 47349 590 47405
rect 646 47349 714 47405
rect 770 47349 838 47405
rect 894 47349 1000 47405
rect 0 47281 1000 47349
rect 0 47225 94 47281
rect 150 47225 218 47281
rect 274 47225 342 47281
rect 398 47225 466 47281
rect 522 47225 590 47281
rect 646 47225 714 47281
rect 770 47225 838 47281
rect 894 47225 1000 47281
rect 0 47157 1000 47225
rect 0 47101 94 47157
rect 150 47101 218 47157
rect 274 47101 342 47157
rect 398 47101 466 47157
rect 522 47101 590 47157
rect 646 47101 714 47157
rect 770 47101 838 47157
rect 894 47101 1000 47157
rect 0 47033 1000 47101
rect 0 46977 94 47033
rect 150 46977 218 47033
rect 274 46977 342 47033
rect 398 46977 466 47033
rect 522 46977 590 47033
rect 646 46977 714 47033
rect 770 46977 838 47033
rect 894 46977 1000 47033
rect 0 46909 1000 46977
rect 0 46853 94 46909
rect 150 46853 218 46909
rect 274 46853 342 46909
rect 398 46853 466 46909
rect 522 46853 590 46909
rect 646 46853 714 46909
rect 770 46853 838 46909
rect 894 46853 1000 46909
rect 0 46785 1000 46853
rect 0 46729 94 46785
rect 150 46729 218 46785
rect 274 46729 342 46785
rect 398 46729 466 46785
rect 522 46729 590 46785
rect 646 46729 714 46785
rect 770 46729 838 46785
rect 894 46729 1000 46785
rect 0 46661 1000 46729
rect 0 46605 94 46661
rect 150 46605 218 46661
rect 274 46605 342 46661
rect 398 46605 466 46661
rect 522 46605 590 46661
rect 646 46605 714 46661
rect 770 46605 838 46661
rect 894 46605 1000 46661
rect 0 46537 1000 46605
rect 0 46481 94 46537
rect 150 46481 218 46537
rect 274 46481 342 46537
rect 398 46481 466 46537
rect 522 46481 590 46537
rect 646 46481 714 46537
rect 770 46481 838 46537
rect 894 46481 1000 46537
rect 0 46413 1000 46481
rect 0 46357 94 46413
rect 150 46357 218 46413
rect 274 46357 342 46413
rect 398 46357 466 46413
rect 522 46357 590 46413
rect 646 46357 714 46413
rect 770 46357 838 46413
rect 894 46357 1000 46413
rect 0 46289 1000 46357
rect 0 46233 94 46289
rect 150 46233 218 46289
rect 274 46233 342 46289
rect 398 46233 466 46289
rect 522 46233 590 46289
rect 646 46233 714 46289
rect 770 46233 838 46289
rect 894 46233 1000 46289
rect 0 46165 1000 46233
rect 0 46109 94 46165
rect 150 46109 218 46165
rect 274 46109 342 46165
rect 398 46109 466 46165
rect 522 46109 590 46165
rect 646 46109 714 46165
rect 770 46109 838 46165
rect 894 46109 1000 46165
rect 0 46099 1000 46109
rect 0 46000 200 46099
rect 800 46000 1000 46099
rect 0 45707 200 45800
rect 800 45707 1000 45800
rect 0 45697 1000 45707
rect 0 45641 94 45697
rect 150 45641 218 45697
rect 274 45641 342 45697
rect 398 45641 466 45697
rect 522 45641 590 45697
rect 646 45641 714 45697
rect 770 45641 838 45697
rect 894 45641 1000 45697
rect 0 45573 1000 45641
rect 0 45517 94 45573
rect 150 45517 218 45573
rect 274 45517 342 45573
rect 398 45517 466 45573
rect 522 45517 590 45573
rect 646 45517 714 45573
rect 770 45517 838 45573
rect 894 45517 1000 45573
rect 0 45449 1000 45517
rect 0 45393 94 45449
rect 150 45393 218 45449
rect 274 45393 342 45449
rect 398 45393 466 45449
rect 522 45393 590 45449
rect 646 45393 714 45449
rect 770 45393 838 45449
rect 894 45393 1000 45449
rect 0 45325 1000 45393
rect 0 45269 94 45325
rect 150 45269 218 45325
rect 274 45269 342 45325
rect 398 45269 466 45325
rect 522 45269 590 45325
rect 646 45269 714 45325
rect 770 45269 838 45325
rect 894 45269 1000 45325
rect 0 45201 1000 45269
rect 0 45145 94 45201
rect 150 45145 218 45201
rect 274 45145 342 45201
rect 398 45145 466 45201
rect 522 45145 590 45201
rect 646 45145 714 45201
rect 770 45145 838 45201
rect 894 45145 1000 45201
rect 0 45077 1000 45145
rect 0 45021 94 45077
rect 150 45021 218 45077
rect 274 45021 342 45077
rect 398 45021 466 45077
rect 522 45021 590 45077
rect 646 45021 714 45077
rect 770 45021 838 45077
rect 894 45021 1000 45077
rect 0 44953 1000 45021
rect 0 44897 94 44953
rect 150 44897 218 44953
rect 274 44897 342 44953
rect 398 44897 466 44953
rect 522 44897 590 44953
rect 646 44897 714 44953
rect 770 44897 838 44953
rect 894 44897 1000 44953
rect 0 44829 1000 44897
rect 0 44773 94 44829
rect 150 44773 218 44829
rect 274 44773 342 44829
rect 398 44773 466 44829
rect 522 44773 590 44829
rect 646 44773 714 44829
rect 770 44773 838 44829
rect 894 44773 1000 44829
rect 0 44705 1000 44773
rect 0 44649 94 44705
rect 150 44649 218 44705
rect 274 44649 342 44705
rect 398 44649 466 44705
rect 522 44649 590 44705
rect 646 44649 714 44705
rect 770 44649 838 44705
rect 894 44649 1000 44705
rect 0 44581 1000 44649
rect 0 44525 94 44581
rect 150 44525 218 44581
rect 274 44525 342 44581
rect 398 44525 466 44581
rect 522 44525 590 44581
rect 646 44525 714 44581
rect 770 44525 838 44581
rect 894 44525 1000 44581
rect 0 44457 1000 44525
rect 0 44401 94 44457
rect 150 44401 218 44457
rect 274 44401 342 44457
rect 398 44401 466 44457
rect 522 44401 590 44457
rect 646 44401 714 44457
rect 770 44401 838 44457
rect 894 44401 1000 44457
rect 0 44333 1000 44401
rect 0 44277 94 44333
rect 150 44277 218 44333
rect 274 44277 342 44333
rect 398 44277 466 44333
rect 522 44277 590 44333
rect 646 44277 714 44333
rect 770 44277 838 44333
rect 894 44277 1000 44333
rect 0 44209 1000 44277
rect 0 44153 94 44209
rect 150 44153 218 44209
rect 274 44153 342 44209
rect 398 44153 466 44209
rect 522 44153 590 44209
rect 646 44153 714 44209
rect 770 44153 838 44209
rect 894 44153 1000 44209
rect 0 44085 1000 44153
rect 0 44029 94 44085
rect 150 44029 218 44085
rect 274 44029 342 44085
rect 398 44029 466 44085
rect 522 44029 590 44085
rect 646 44029 714 44085
rect 770 44029 838 44085
rect 894 44029 1000 44085
rect 0 43961 1000 44029
rect 0 43905 94 43961
rect 150 43905 218 43961
rect 274 43905 342 43961
rect 398 43905 466 43961
rect 522 43905 590 43961
rect 646 43905 714 43961
rect 770 43905 838 43961
rect 894 43905 1000 43961
rect 0 43837 1000 43905
rect 0 43781 94 43837
rect 150 43781 218 43837
rect 274 43781 342 43837
rect 398 43781 466 43837
rect 522 43781 590 43837
rect 646 43781 714 43837
rect 770 43781 838 43837
rect 894 43781 1000 43837
rect 0 43713 1000 43781
rect 0 43657 94 43713
rect 150 43657 218 43713
rect 274 43657 342 43713
rect 398 43657 466 43713
rect 522 43657 590 43713
rect 646 43657 714 43713
rect 770 43657 838 43713
rect 894 43657 1000 43713
rect 0 43589 1000 43657
rect 0 43533 94 43589
rect 150 43533 218 43589
rect 274 43533 342 43589
rect 398 43533 466 43589
rect 522 43533 590 43589
rect 646 43533 714 43589
rect 770 43533 838 43589
rect 894 43533 1000 43589
rect 0 43465 1000 43533
rect 0 43409 94 43465
rect 150 43409 218 43465
rect 274 43409 342 43465
rect 398 43409 466 43465
rect 522 43409 590 43465
rect 646 43409 714 43465
rect 770 43409 838 43465
rect 894 43409 1000 43465
rect 0 43341 1000 43409
rect 0 43285 94 43341
rect 150 43285 218 43341
rect 274 43285 342 43341
rect 398 43285 466 43341
rect 522 43285 590 43341
rect 646 43285 714 43341
rect 770 43285 838 43341
rect 894 43285 1000 43341
rect 0 43217 1000 43285
rect 0 43161 94 43217
rect 150 43161 218 43217
rect 274 43161 342 43217
rect 398 43161 466 43217
rect 522 43161 590 43217
rect 646 43161 714 43217
rect 770 43161 838 43217
rect 894 43161 1000 43217
rect 0 43093 1000 43161
rect 0 43037 94 43093
rect 150 43037 218 43093
rect 274 43037 342 43093
rect 398 43037 466 43093
rect 522 43037 590 43093
rect 646 43037 714 43093
rect 770 43037 838 43093
rect 894 43037 1000 43093
rect 0 42969 1000 43037
rect 0 42913 94 42969
rect 150 42913 218 42969
rect 274 42913 342 42969
rect 398 42913 466 42969
rect 522 42913 590 42969
rect 646 42913 714 42969
rect 770 42913 838 42969
rect 894 42913 1000 42969
rect 0 42903 1000 42913
rect 0 42800 200 42903
rect 800 42800 1000 42903
rect 0 42494 200 42600
rect 800 42494 1000 42600
rect 0 42484 1000 42494
rect 0 42428 95 42484
rect 151 42428 219 42484
rect 275 42428 343 42484
rect 399 42428 467 42484
rect 523 42428 591 42484
rect 647 42428 715 42484
rect 771 42428 839 42484
rect 895 42428 1000 42484
rect 0 42360 1000 42428
rect 0 42304 95 42360
rect 151 42304 219 42360
rect 275 42304 343 42360
rect 399 42304 467 42360
rect 523 42304 591 42360
rect 647 42304 715 42360
rect 771 42304 839 42360
rect 895 42304 1000 42360
rect 0 42236 1000 42304
rect 0 42180 95 42236
rect 151 42180 219 42236
rect 275 42180 343 42236
rect 399 42180 467 42236
rect 523 42180 591 42236
rect 647 42180 715 42236
rect 771 42180 839 42236
rect 895 42180 1000 42236
rect 0 42112 1000 42180
rect 0 42056 95 42112
rect 151 42056 219 42112
rect 275 42056 343 42112
rect 399 42056 467 42112
rect 523 42056 591 42112
rect 647 42056 715 42112
rect 771 42056 839 42112
rect 895 42056 1000 42112
rect 0 41988 1000 42056
rect 0 41932 95 41988
rect 151 41932 219 41988
rect 275 41932 343 41988
rect 399 41932 467 41988
rect 523 41932 591 41988
rect 647 41932 715 41988
rect 771 41932 839 41988
rect 895 41932 1000 41988
rect 0 41864 1000 41932
rect 0 41808 95 41864
rect 151 41808 219 41864
rect 275 41808 343 41864
rect 399 41808 467 41864
rect 523 41808 591 41864
rect 647 41808 715 41864
rect 771 41808 839 41864
rect 895 41808 1000 41864
rect 0 41740 1000 41808
rect 0 41684 95 41740
rect 151 41684 219 41740
rect 275 41684 343 41740
rect 399 41684 467 41740
rect 523 41684 591 41740
rect 647 41684 715 41740
rect 771 41684 839 41740
rect 895 41684 1000 41740
rect 0 41616 1000 41684
rect 0 41560 95 41616
rect 151 41560 219 41616
rect 275 41560 343 41616
rect 399 41560 467 41616
rect 523 41560 591 41616
rect 647 41560 715 41616
rect 771 41560 839 41616
rect 895 41560 1000 41616
rect 0 41492 1000 41560
rect 0 41436 95 41492
rect 151 41436 219 41492
rect 275 41436 343 41492
rect 399 41436 467 41492
rect 523 41436 591 41492
rect 647 41436 715 41492
rect 771 41436 839 41492
rect 895 41436 1000 41492
rect 0 41368 1000 41436
rect 0 41312 95 41368
rect 151 41312 219 41368
rect 275 41312 343 41368
rect 399 41312 467 41368
rect 523 41312 591 41368
rect 647 41312 715 41368
rect 771 41312 839 41368
rect 895 41312 1000 41368
rect 0 41302 1000 41312
rect 0 41200 200 41302
rect 800 41200 1000 41302
rect 0 40906 200 41000
rect 800 40906 1000 41000
rect 0 40896 1000 40906
rect 0 40840 95 40896
rect 151 40840 219 40896
rect 275 40840 343 40896
rect 399 40840 467 40896
rect 523 40840 591 40896
rect 647 40840 715 40896
rect 771 40840 839 40896
rect 895 40840 1000 40896
rect 0 40772 1000 40840
rect 0 40716 95 40772
rect 151 40716 219 40772
rect 275 40716 343 40772
rect 399 40716 467 40772
rect 523 40716 591 40772
rect 647 40716 715 40772
rect 771 40716 839 40772
rect 895 40716 1000 40772
rect 0 40648 1000 40716
rect 0 40592 95 40648
rect 151 40592 219 40648
rect 275 40592 343 40648
rect 399 40592 467 40648
rect 523 40592 591 40648
rect 647 40592 715 40648
rect 771 40592 839 40648
rect 895 40592 1000 40648
rect 0 40524 1000 40592
rect 0 40468 95 40524
rect 151 40468 219 40524
rect 275 40468 343 40524
rect 399 40468 467 40524
rect 523 40468 591 40524
rect 647 40468 715 40524
rect 771 40468 839 40524
rect 895 40468 1000 40524
rect 0 40400 1000 40468
rect 0 40344 95 40400
rect 151 40344 219 40400
rect 275 40344 343 40400
rect 399 40344 467 40400
rect 523 40344 591 40400
rect 647 40344 715 40400
rect 771 40344 839 40400
rect 895 40344 1000 40400
rect 0 40276 1000 40344
rect 0 40220 95 40276
rect 151 40220 219 40276
rect 275 40220 343 40276
rect 399 40220 467 40276
rect 523 40220 591 40276
rect 647 40220 715 40276
rect 771 40220 839 40276
rect 895 40220 1000 40276
rect 0 40152 1000 40220
rect 0 40096 95 40152
rect 151 40096 219 40152
rect 275 40096 343 40152
rect 399 40096 467 40152
rect 523 40096 591 40152
rect 647 40096 715 40152
rect 771 40096 839 40152
rect 895 40096 1000 40152
rect 0 40028 1000 40096
rect 0 39972 95 40028
rect 151 39972 219 40028
rect 275 39972 343 40028
rect 399 39972 467 40028
rect 523 39972 591 40028
rect 647 39972 715 40028
rect 771 39972 839 40028
rect 895 39972 1000 40028
rect 0 39904 1000 39972
rect 0 39848 95 39904
rect 151 39848 219 39904
rect 275 39848 343 39904
rect 399 39848 467 39904
rect 523 39848 591 39904
rect 647 39848 715 39904
rect 771 39848 839 39904
rect 895 39848 1000 39904
rect 0 39780 1000 39848
rect 0 39724 95 39780
rect 151 39724 219 39780
rect 275 39724 343 39780
rect 399 39724 467 39780
rect 523 39724 591 39780
rect 647 39724 715 39780
rect 771 39724 839 39780
rect 895 39724 1000 39780
rect 0 39714 1000 39724
rect 0 39600 200 39714
rect 800 39600 1000 39714
rect 0 39314 200 39400
rect 800 39314 1000 39400
rect 0 39304 1000 39314
rect 0 39248 94 39304
rect 150 39248 218 39304
rect 274 39248 342 39304
rect 398 39248 466 39304
rect 522 39248 590 39304
rect 646 39248 714 39304
rect 770 39248 838 39304
rect 894 39248 1000 39304
rect 0 39180 1000 39248
rect 0 39124 94 39180
rect 150 39124 218 39180
rect 274 39124 342 39180
rect 398 39124 466 39180
rect 522 39124 590 39180
rect 646 39124 714 39180
rect 770 39124 838 39180
rect 894 39124 1000 39180
rect 0 39056 1000 39124
rect 0 39000 94 39056
rect 150 39000 218 39056
rect 274 39000 342 39056
rect 398 39000 466 39056
rect 522 39000 590 39056
rect 646 39000 714 39056
rect 770 39000 838 39056
rect 894 39000 1000 39056
rect 0 38932 1000 39000
rect 0 38876 94 38932
rect 150 38876 218 38932
rect 274 38876 342 38932
rect 398 38876 466 38932
rect 522 38876 590 38932
rect 646 38876 714 38932
rect 770 38876 838 38932
rect 894 38876 1000 38932
rect 0 38808 1000 38876
rect 0 38752 94 38808
rect 150 38752 218 38808
rect 274 38752 342 38808
rect 398 38752 466 38808
rect 522 38752 590 38808
rect 646 38752 714 38808
rect 770 38752 838 38808
rect 894 38752 1000 38808
rect 0 38684 1000 38752
rect 0 38628 94 38684
rect 150 38628 218 38684
rect 274 38628 342 38684
rect 398 38628 466 38684
rect 522 38628 590 38684
rect 646 38628 714 38684
rect 770 38628 838 38684
rect 894 38628 1000 38684
rect 0 38560 1000 38628
rect 0 38504 94 38560
rect 150 38504 218 38560
rect 274 38504 342 38560
rect 398 38504 466 38560
rect 522 38504 590 38560
rect 646 38504 714 38560
rect 770 38504 838 38560
rect 894 38504 1000 38560
rect 0 38436 1000 38504
rect 0 38380 94 38436
rect 150 38380 218 38436
rect 274 38380 342 38436
rect 398 38380 466 38436
rect 522 38380 590 38436
rect 646 38380 714 38436
rect 770 38380 838 38436
rect 894 38380 1000 38436
rect 0 38312 1000 38380
rect 0 38256 94 38312
rect 150 38256 218 38312
rect 274 38256 342 38312
rect 398 38256 466 38312
rect 522 38256 590 38312
rect 646 38256 714 38312
rect 770 38256 838 38312
rect 894 38256 1000 38312
rect 0 38188 1000 38256
rect 0 38132 94 38188
rect 150 38132 218 38188
rect 274 38132 342 38188
rect 398 38132 466 38188
rect 522 38132 590 38188
rect 646 38132 714 38188
rect 770 38132 838 38188
rect 894 38132 1000 38188
rect 0 38064 1000 38132
rect 0 38008 94 38064
rect 150 38008 218 38064
rect 274 38008 342 38064
rect 398 38008 466 38064
rect 522 38008 590 38064
rect 646 38008 714 38064
rect 770 38008 838 38064
rect 894 38008 1000 38064
rect 0 37940 1000 38008
rect 0 37884 94 37940
rect 150 37884 218 37940
rect 274 37884 342 37940
rect 398 37884 466 37940
rect 522 37884 590 37940
rect 646 37884 714 37940
rect 770 37884 838 37940
rect 894 37884 1000 37940
rect 0 37816 1000 37884
rect 0 37760 94 37816
rect 150 37760 218 37816
rect 274 37760 342 37816
rect 398 37760 466 37816
rect 522 37760 590 37816
rect 646 37760 714 37816
rect 770 37760 838 37816
rect 894 37760 1000 37816
rect 0 37692 1000 37760
rect 0 37636 94 37692
rect 150 37636 218 37692
rect 274 37636 342 37692
rect 398 37636 466 37692
rect 522 37636 590 37692
rect 646 37636 714 37692
rect 770 37636 838 37692
rect 894 37636 1000 37692
rect 0 37568 1000 37636
rect 0 37512 94 37568
rect 150 37512 218 37568
rect 274 37512 342 37568
rect 398 37512 466 37568
rect 522 37512 590 37568
rect 646 37512 714 37568
rect 770 37512 838 37568
rect 894 37512 1000 37568
rect 0 37444 1000 37512
rect 0 37388 94 37444
rect 150 37388 218 37444
rect 274 37388 342 37444
rect 398 37388 466 37444
rect 522 37388 590 37444
rect 646 37388 714 37444
rect 770 37388 838 37444
rect 894 37388 1000 37444
rect 0 37320 1000 37388
rect 0 37264 94 37320
rect 150 37264 218 37320
rect 274 37264 342 37320
rect 398 37264 466 37320
rect 522 37264 590 37320
rect 646 37264 714 37320
rect 770 37264 838 37320
rect 894 37264 1000 37320
rect 0 37196 1000 37264
rect 0 37140 94 37196
rect 150 37140 218 37196
rect 274 37140 342 37196
rect 398 37140 466 37196
rect 522 37140 590 37196
rect 646 37140 714 37196
rect 770 37140 838 37196
rect 894 37140 1000 37196
rect 0 37072 1000 37140
rect 0 37016 94 37072
rect 150 37016 218 37072
rect 274 37016 342 37072
rect 398 37016 466 37072
rect 522 37016 590 37072
rect 646 37016 714 37072
rect 770 37016 838 37072
rect 894 37016 1000 37072
rect 0 36948 1000 37016
rect 0 36892 94 36948
rect 150 36892 218 36948
rect 274 36892 342 36948
rect 398 36892 466 36948
rect 522 36892 590 36948
rect 646 36892 714 36948
rect 770 36892 838 36948
rect 894 36892 1000 36948
rect 0 36824 1000 36892
rect 0 36768 94 36824
rect 150 36768 218 36824
rect 274 36768 342 36824
rect 398 36768 466 36824
rect 522 36768 590 36824
rect 646 36768 714 36824
rect 770 36768 838 36824
rect 894 36768 1000 36824
rect 0 36700 1000 36768
rect 0 36644 94 36700
rect 150 36644 218 36700
rect 274 36644 342 36700
rect 398 36644 466 36700
rect 522 36644 590 36700
rect 646 36644 714 36700
rect 770 36644 838 36700
rect 894 36644 1000 36700
rect 0 36576 1000 36644
rect 0 36520 94 36576
rect 150 36520 218 36576
rect 274 36520 342 36576
rect 398 36520 466 36576
rect 522 36520 590 36576
rect 646 36520 714 36576
rect 770 36520 838 36576
rect 894 36520 1000 36576
rect 0 36510 1000 36520
rect 0 36400 200 36510
rect 800 36400 1000 36510
rect 0 36104 200 36200
rect 800 36104 1000 36200
rect 0 36094 1000 36104
rect 0 36038 94 36094
rect 150 36038 218 36094
rect 274 36038 342 36094
rect 398 36038 466 36094
rect 522 36038 590 36094
rect 646 36038 714 36094
rect 770 36038 838 36094
rect 894 36038 1000 36094
rect 0 35970 1000 36038
rect 0 35914 94 35970
rect 150 35914 218 35970
rect 274 35914 342 35970
rect 398 35914 466 35970
rect 522 35914 590 35970
rect 646 35914 714 35970
rect 770 35914 838 35970
rect 894 35914 1000 35970
rect 0 35846 1000 35914
rect 0 35790 94 35846
rect 150 35790 218 35846
rect 274 35790 342 35846
rect 398 35790 466 35846
rect 522 35790 590 35846
rect 646 35790 714 35846
rect 770 35790 838 35846
rect 894 35790 1000 35846
rect 0 35722 1000 35790
rect 0 35666 94 35722
rect 150 35666 218 35722
rect 274 35666 342 35722
rect 398 35666 466 35722
rect 522 35666 590 35722
rect 646 35666 714 35722
rect 770 35666 838 35722
rect 894 35666 1000 35722
rect 0 35598 1000 35666
rect 0 35542 94 35598
rect 150 35542 218 35598
rect 274 35542 342 35598
rect 398 35542 466 35598
rect 522 35542 590 35598
rect 646 35542 714 35598
rect 770 35542 838 35598
rect 894 35542 1000 35598
rect 0 35474 1000 35542
rect 0 35418 94 35474
rect 150 35418 218 35474
rect 274 35418 342 35474
rect 398 35418 466 35474
rect 522 35418 590 35474
rect 646 35418 714 35474
rect 770 35418 838 35474
rect 894 35418 1000 35474
rect 0 35350 1000 35418
rect 0 35294 94 35350
rect 150 35294 218 35350
rect 274 35294 342 35350
rect 398 35294 466 35350
rect 522 35294 590 35350
rect 646 35294 714 35350
rect 770 35294 838 35350
rect 894 35294 1000 35350
rect 0 35226 1000 35294
rect 0 35170 94 35226
rect 150 35170 218 35226
rect 274 35170 342 35226
rect 398 35170 466 35226
rect 522 35170 590 35226
rect 646 35170 714 35226
rect 770 35170 838 35226
rect 894 35170 1000 35226
rect 0 35102 1000 35170
rect 0 35046 94 35102
rect 150 35046 218 35102
rect 274 35046 342 35102
rect 398 35046 466 35102
rect 522 35046 590 35102
rect 646 35046 714 35102
rect 770 35046 838 35102
rect 894 35046 1000 35102
rect 0 34978 1000 35046
rect 0 34922 94 34978
rect 150 34922 218 34978
rect 274 34922 342 34978
rect 398 34922 466 34978
rect 522 34922 590 34978
rect 646 34922 714 34978
rect 770 34922 838 34978
rect 894 34922 1000 34978
rect 0 34854 1000 34922
rect 0 34798 94 34854
rect 150 34798 218 34854
rect 274 34798 342 34854
rect 398 34798 466 34854
rect 522 34798 590 34854
rect 646 34798 714 34854
rect 770 34798 838 34854
rect 894 34798 1000 34854
rect 0 34730 1000 34798
rect 0 34674 94 34730
rect 150 34674 218 34730
rect 274 34674 342 34730
rect 398 34674 466 34730
rect 522 34674 590 34730
rect 646 34674 714 34730
rect 770 34674 838 34730
rect 894 34674 1000 34730
rect 0 34606 1000 34674
rect 0 34550 94 34606
rect 150 34550 218 34606
rect 274 34550 342 34606
rect 398 34550 466 34606
rect 522 34550 590 34606
rect 646 34550 714 34606
rect 770 34550 838 34606
rect 894 34550 1000 34606
rect 0 34482 1000 34550
rect 0 34426 94 34482
rect 150 34426 218 34482
rect 274 34426 342 34482
rect 398 34426 466 34482
rect 522 34426 590 34482
rect 646 34426 714 34482
rect 770 34426 838 34482
rect 894 34426 1000 34482
rect 0 34358 1000 34426
rect 0 34302 94 34358
rect 150 34302 218 34358
rect 274 34302 342 34358
rect 398 34302 466 34358
rect 522 34302 590 34358
rect 646 34302 714 34358
rect 770 34302 838 34358
rect 894 34302 1000 34358
rect 0 34234 1000 34302
rect 0 34178 94 34234
rect 150 34178 218 34234
rect 274 34178 342 34234
rect 398 34178 466 34234
rect 522 34178 590 34234
rect 646 34178 714 34234
rect 770 34178 838 34234
rect 894 34178 1000 34234
rect 0 34110 1000 34178
rect 0 34054 94 34110
rect 150 34054 218 34110
rect 274 34054 342 34110
rect 398 34054 466 34110
rect 522 34054 590 34110
rect 646 34054 714 34110
rect 770 34054 838 34110
rect 894 34054 1000 34110
rect 0 33986 1000 34054
rect 0 33930 94 33986
rect 150 33930 218 33986
rect 274 33930 342 33986
rect 398 33930 466 33986
rect 522 33930 590 33986
rect 646 33930 714 33986
rect 770 33930 838 33986
rect 894 33930 1000 33986
rect 0 33862 1000 33930
rect 0 33806 94 33862
rect 150 33806 218 33862
rect 274 33806 342 33862
rect 398 33806 466 33862
rect 522 33806 590 33862
rect 646 33806 714 33862
rect 770 33806 838 33862
rect 894 33806 1000 33862
rect 0 33738 1000 33806
rect 0 33682 94 33738
rect 150 33682 218 33738
rect 274 33682 342 33738
rect 398 33682 466 33738
rect 522 33682 590 33738
rect 646 33682 714 33738
rect 770 33682 838 33738
rect 894 33682 1000 33738
rect 0 33614 1000 33682
rect 0 33558 94 33614
rect 150 33558 218 33614
rect 274 33558 342 33614
rect 398 33558 466 33614
rect 522 33558 590 33614
rect 646 33558 714 33614
rect 770 33558 838 33614
rect 894 33558 1000 33614
rect 0 33490 1000 33558
rect 0 33434 94 33490
rect 150 33434 218 33490
rect 274 33434 342 33490
rect 398 33434 466 33490
rect 522 33434 590 33490
rect 646 33434 714 33490
rect 770 33434 838 33490
rect 894 33434 1000 33490
rect 0 33366 1000 33434
rect 0 33310 94 33366
rect 150 33310 218 33366
rect 274 33310 342 33366
rect 398 33310 466 33366
rect 522 33310 590 33366
rect 646 33310 714 33366
rect 770 33310 838 33366
rect 894 33310 1000 33366
rect 0 33300 1000 33310
rect 0 33200 200 33300
rect 800 33200 1000 33300
rect 0 32912 200 33000
rect 800 32912 1000 33000
rect 0 32902 1000 32912
rect 0 32846 94 32902
rect 150 32846 218 32902
rect 274 32846 342 32902
rect 398 32846 466 32902
rect 522 32846 590 32902
rect 646 32846 714 32902
rect 770 32846 838 32902
rect 894 32846 1000 32902
rect 0 32778 1000 32846
rect 0 32722 94 32778
rect 150 32722 218 32778
rect 274 32722 342 32778
rect 398 32722 466 32778
rect 522 32722 590 32778
rect 646 32722 714 32778
rect 770 32722 838 32778
rect 894 32722 1000 32778
rect 0 32654 1000 32722
rect 0 32598 94 32654
rect 150 32598 218 32654
rect 274 32598 342 32654
rect 398 32598 466 32654
rect 522 32598 590 32654
rect 646 32598 714 32654
rect 770 32598 838 32654
rect 894 32598 1000 32654
rect 0 32530 1000 32598
rect 0 32474 94 32530
rect 150 32474 218 32530
rect 274 32474 342 32530
rect 398 32474 466 32530
rect 522 32474 590 32530
rect 646 32474 714 32530
rect 770 32474 838 32530
rect 894 32474 1000 32530
rect 0 32406 1000 32474
rect 0 32350 94 32406
rect 150 32350 218 32406
rect 274 32350 342 32406
rect 398 32350 466 32406
rect 522 32350 590 32406
rect 646 32350 714 32406
rect 770 32350 838 32406
rect 894 32350 1000 32406
rect 0 32282 1000 32350
rect 0 32226 94 32282
rect 150 32226 218 32282
rect 274 32226 342 32282
rect 398 32226 466 32282
rect 522 32226 590 32282
rect 646 32226 714 32282
rect 770 32226 838 32282
rect 894 32226 1000 32282
rect 0 32158 1000 32226
rect 0 32102 94 32158
rect 150 32102 218 32158
rect 274 32102 342 32158
rect 398 32102 466 32158
rect 522 32102 590 32158
rect 646 32102 714 32158
rect 770 32102 838 32158
rect 894 32102 1000 32158
rect 0 32034 1000 32102
rect 0 31978 94 32034
rect 150 31978 218 32034
rect 274 31978 342 32034
rect 398 31978 466 32034
rect 522 31978 590 32034
rect 646 31978 714 32034
rect 770 31978 838 32034
rect 894 31978 1000 32034
rect 0 31910 1000 31978
rect 0 31854 94 31910
rect 150 31854 218 31910
rect 274 31854 342 31910
rect 398 31854 466 31910
rect 522 31854 590 31910
rect 646 31854 714 31910
rect 770 31854 838 31910
rect 894 31854 1000 31910
rect 0 31786 1000 31854
rect 0 31730 94 31786
rect 150 31730 218 31786
rect 274 31730 342 31786
rect 398 31730 466 31786
rect 522 31730 590 31786
rect 646 31730 714 31786
rect 770 31730 838 31786
rect 894 31730 1000 31786
rect 0 31662 1000 31730
rect 0 31606 94 31662
rect 150 31606 218 31662
rect 274 31606 342 31662
rect 398 31606 466 31662
rect 522 31606 590 31662
rect 646 31606 714 31662
rect 770 31606 838 31662
rect 894 31606 1000 31662
rect 0 31538 1000 31606
rect 0 31482 94 31538
rect 150 31482 218 31538
rect 274 31482 342 31538
rect 398 31482 466 31538
rect 522 31482 590 31538
rect 646 31482 714 31538
rect 770 31482 838 31538
rect 894 31482 1000 31538
rect 0 31414 1000 31482
rect 0 31358 94 31414
rect 150 31358 218 31414
rect 274 31358 342 31414
rect 398 31358 466 31414
rect 522 31358 590 31414
rect 646 31358 714 31414
rect 770 31358 838 31414
rect 894 31358 1000 31414
rect 0 31290 1000 31358
rect 0 31234 94 31290
rect 150 31234 218 31290
rect 274 31234 342 31290
rect 398 31234 466 31290
rect 522 31234 590 31290
rect 646 31234 714 31290
rect 770 31234 838 31290
rect 894 31234 1000 31290
rect 0 31166 1000 31234
rect 0 31110 94 31166
rect 150 31110 218 31166
rect 274 31110 342 31166
rect 398 31110 466 31166
rect 522 31110 590 31166
rect 646 31110 714 31166
rect 770 31110 838 31166
rect 894 31110 1000 31166
rect 0 31042 1000 31110
rect 0 30986 94 31042
rect 150 30986 218 31042
rect 274 30986 342 31042
rect 398 30986 466 31042
rect 522 30986 590 31042
rect 646 30986 714 31042
rect 770 30986 838 31042
rect 894 30986 1000 31042
rect 0 30918 1000 30986
rect 0 30862 94 30918
rect 150 30862 218 30918
rect 274 30862 342 30918
rect 398 30862 466 30918
rect 522 30862 590 30918
rect 646 30862 714 30918
rect 770 30862 838 30918
rect 894 30862 1000 30918
rect 0 30794 1000 30862
rect 0 30738 94 30794
rect 150 30738 218 30794
rect 274 30738 342 30794
rect 398 30738 466 30794
rect 522 30738 590 30794
rect 646 30738 714 30794
rect 770 30738 838 30794
rect 894 30738 1000 30794
rect 0 30670 1000 30738
rect 0 30614 94 30670
rect 150 30614 218 30670
rect 274 30614 342 30670
rect 398 30614 466 30670
rect 522 30614 590 30670
rect 646 30614 714 30670
rect 770 30614 838 30670
rect 894 30614 1000 30670
rect 0 30546 1000 30614
rect 0 30490 94 30546
rect 150 30490 218 30546
rect 274 30490 342 30546
rect 398 30490 466 30546
rect 522 30490 590 30546
rect 646 30490 714 30546
rect 770 30490 838 30546
rect 894 30490 1000 30546
rect 0 30422 1000 30490
rect 0 30366 94 30422
rect 150 30366 218 30422
rect 274 30366 342 30422
rect 398 30366 466 30422
rect 522 30366 590 30422
rect 646 30366 714 30422
rect 770 30366 838 30422
rect 894 30366 1000 30422
rect 0 30298 1000 30366
rect 0 30242 94 30298
rect 150 30242 218 30298
rect 274 30242 342 30298
rect 398 30242 466 30298
rect 522 30242 590 30298
rect 646 30242 714 30298
rect 770 30242 838 30298
rect 894 30242 1000 30298
rect 0 30174 1000 30242
rect 0 30118 94 30174
rect 150 30118 218 30174
rect 274 30118 342 30174
rect 398 30118 466 30174
rect 522 30118 590 30174
rect 646 30118 714 30174
rect 770 30118 838 30174
rect 894 30118 1000 30174
rect 0 30108 1000 30118
rect 0 30000 200 30108
rect 800 30000 1000 30108
rect 0 29695 200 29800
rect 800 29695 1000 29800
rect 0 29685 1000 29695
rect 0 29629 94 29685
rect 150 29629 218 29685
rect 274 29629 342 29685
rect 398 29629 466 29685
rect 522 29629 590 29685
rect 646 29629 714 29685
rect 770 29629 838 29685
rect 894 29629 1000 29685
rect 0 29561 1000 29629
rect 0 29505 94 29561
rect 150 29505 218 29561
rect 274 29505 342 29561
rect 398 29505 466 29561
rect 522 29505 590 29561
rect 646 29505 714 29561
rect 770 29505 838 29561
rect 894 29505 1000 29561
rect 0 29437 1000 29505
rect 0 29381 94 29437
rect 150 29381 218 29437
rect 274 29381 342 29437
rect 398 29381 466 29437
rect 522 29381 590 29437
rect 646 29381 714 29437
rect 770 29381 838 29437
rect 894 29381 1000 29437
rect 0 29313 1000 29381
rect 0 29257 94 29313
rect 150 29257 218 29313
rect 274 29257 342 29313
rect 398 29257 466 29313
rect 522 29257 590 29313
rect 646 29257 714 29313
rect 770 29257 838 29313
rect 894 29257 1000 29313
rect 0 29189 1000 29257
rect 0 29133 94 29189
rect 150 29133 218 29189
rect 274 29133 342 29189
rect 398 29133 466 29189
rect 522 29133 590 29189
rect 646 29133 714 29189
rect 770 29133 838 29189
rect 894 29133 1000 29189
rect 0 29065 1000 29133
rect 0 29009 94 29065
rect 150 29009 218 29065
rect 274 29009 342 29065
rect 398 29009 466 29065
rect 522 29009 590 29065
rect 646 29009 714 29065
rect 770 29009 838 29065
rect 894 29009 1000 29065
rect 0 28941 1000 29009
rect 0 28885 94 28941
rect 150 28885 218 28941
rect 274 28885 342 28941
rect 398 28885 466 28941
rect 522 28885 590 28941
rect 646 28885 714 28941
rect 770 28885 838 28941
rect 894 28885 1000 28941
rect 0 28817 1000 28885
rect 0 28761 94 28817
rect 150 28761 218 28817
rect 274 28761 342 28817
rect 398 28761 466 28817
rect 522 28761 590 28817
rect 646 28761 714 28817
rect 770 28761 838 28817
rect 894 28761 1000 28817
rect 0 28693 1000 28761
rect 0 28637 94 28693
rect 150 28637 218 28693
rect 274 28637 342 28693
rect 398 28637 466 28693
rect 522 28637 590 28693
rect 646 28637 714 28693
rect 770 28637 838 28693
rect 894 28637 1000 28693
rect 0 28569 1000 28637
rect 0 28513 94 28569
rect 150 28513 218 28569
rect 274 28513 342 28569
rect 398 28513 466 28569
rect 522 28513 590 28569
rect 646 28513 714 28569
rect 770 28513 838 28569
rect 894 28513 1000 28569
rect 0 28445 1000 28513
rect 0 28389 94 28445
rect 150 28389 218 28445
rect 274 28389 342 28445
rect 398 28389 466 28445
rect 522 28389 590 28445
rect 646 28389 714 28445
rect 770 28389 838 28445
rect 894 28389 1000 28445
rect 0 28321 1000 28389
rect 0 28265 94 28321
rect 150 28265 218 28321
rect 274 28265 342 28321
rect 398 28265 466 28321
rect 522 28265 590 28321
rect 646 28265 714 28321
rect 770 28265 838 28321
rect 894 28265 1000 28321
rect 0 28197 1000 28265
rect 0 28141 94 28197
rect 150 28141 218 28197
rect 274 28141 342 28197
rect 398 28141 466 28197
rect 522 28141 590 28197
rect 646 28141 714 28197
rect 770 28141 838 28197
rect 894 28141 1000 28197
rect 0 28073 1000 28141
rect 0 28017 94 28073
rect 150 28017 218 28073
rect 274 28017 342 28073
rect 398 28017 466 28073
rect 522 28017 590 28073
rect 646 28017 714 28073
rect 770 28017 838 28073
rect 894 28017 1000 28073
rect 0 27949 1000 28017
rect 0 27893 94 27949
rect 150 27893 218 27949
rect 274 27893 342 27949
rect 398 27893 466 27949
rect 522 27893 590 27949
rect 646 27893 714 27949
rect 770 27893 838 27949
rect 894 27893 1000 27949
rect 0 27825 1000 27893
rect 0 27769 94 27825
rect 150 27769 218 27825
rect 274 27769 342 27825
rect 398 27769 466 27825
rect 522 27769 590 27825
rect 646 27769 714 27825
rect 770 27769 838 27825
rect 894 27769 1000 27825
rect 0 27701 1000 27769
rect 0 27645 94 27701
rect 150 27645 218 27701
rect 274 27645 342 27701
rect 398 27645 466 27701
rect 522 27645 590 27701
rect 646 27645 714 27701
rect 770 27645 838 27701
rect 894 27645 1000 27701
rect 0 27577 1000 27645
rect 0 27521 94 27577
rect 150 27521 218 27577
rect 274 27521 342 27577
rect 398 27521 466 27577
rect 522 27521 590 27577
rect 646 27521 714 27577
rect 770 27521 838 27577
rect 894 27521 1000 27577
rect 0 27453 1000 27521
rect 0 27397 94 27453
rect 150 27397 218 27453
rect 274 27397 342 27453
rect 398 27397 466 27453
rect 522 27397 590 27453
rect 646 27397 714 27453
rect 770 27397 838 27453
rect 894 27397 1000 27453
rect 0 27329 1000 27397
rect 0 27273 94 27329
rect 150 27273 218 27329
rect 274 27273 342 27329
rect 398 27273 466 27329
rect 522 27273 590 27329
rect 646 27273 714 27329
rect 770 27273 838 27329
rect 894 27273 1000 27329
rect 0 27205 1000 27273
rect 0 27149 94 27205
rect 150 27149 218 27205
rect 274 27149 342 27205
rect 398 27149 466 27205
rect 522 27149 590 27205
rect 646 27149 714 27205
rect 770 27149 838 27205
rect 894 27149 1000 27205
rect 0 27081 1000 27149
rect 0 27025 94 27081
rect 150 27025 218 27081
rect 274 27025 342 27081
rect 398 27025 466 27081
rect 522 27025 590 27081
rect 646 27025 714 27081
rect 770 27025 838 27081
rect 894 27025 1000 27081
rect 0 26957 1000 27025
rect 0 26901 94 26957
rect 150 26901 218 26957
rect 274 26901 342 26957
rect 398 26901 466 26957
rect 522 26901 590 26957
rect 646 26901 714 26957
rect 770 26901 838 26957
rect 894 26901 1000 26957
rect 0 26891 1000 26901
rect 0 26800 200 26891
rect 800 26800 1000 26891
rect 0 26506 200 26600
rect 800 26506 1000 26600
rect 0 26496 1000 26506
rect 0 26440 95 26496
rect 151 26440 219 26496
rect 275 26440 343 26496
rect 399 26440 467 26496
rect 523 26440 591 26496
rect 647 26440 715 26496
rect 771 26440 839 26496
rect 895 26440 1000 26496
rect 0 26372 1000 26440
rect 0 26316 95 26372
rect 151 26316 219 26372
rect 275 26316 343 26372
rect 399 26316 467 26372
rect 523 26316 591 26372
rect 647 26316 715 26372
rect 771 26316 839 26372
rect 895 26316 1000 26372
rect 0 26248 1000 26316
rect 0 26192 95 26248
rect 151 26192 219 26248
rect 275 26192 343 26248
rect 399 26192 467 26248
rect 523 26192 591 26248
rect 647 26192 715 26248
rect 771 26192 839 26248
rect 895 26192 1000 26248
rect 0 26124 1000 26192
rect 0 26068 95 26124
rect 151 26068 219 26124
rect 275 26068 343 26124
rect 399 26068 467 26124
rect 523 26068 591 26124
rect 647 26068 715 26124
rect 771 26068 839 26124
rect 895 26068 1000 26124
rect 0 26000 1000 26068
rect 0 25944 95 26000
rect 151 25944 219 26000
rect 275 25944 343 26000
rect 399 25944 467 26000
rect 523 25944 591 26000
rect 647 25944 715 26000
rect 771 25944 839 26000
rect 895 25944 1000 26000
rect 0 25876 1000 25944
rect 0 25820 95 25876
rect 151 25820 219 25876
rect 275 25820 343 25876
rect 399 25820 467 25876
rect 523 25820 591 25876
rect 647 25820 715 25876
rect 771 25820 839 25876
rect 895 25820 1000 25876
rect 0 25752 1000 25820
rect 0 25696 95 25752
rect 151 25696 219 25752
rect 275 25696 343 25752
rect 399 25696 467 25752
rect 523 25696 591 25752
rect 647 25696 715 25752
rect 771 25696 839 25752
rect 895 25696 1000 25752
rect 0 25628 1000 25696
rect 0 25572 95 25628
rect 151 25572 219 25628
rect 275 25572 343 25628
rect 399 25572 467 25628
rect 523 25572 591 25628
rect 647 25572 715 25628
rect 771 25572 839 25628
rect 895 25572 1000 25628
rect 0 25504 1000 25572
rect 0 25448 95 25504
rect 151 25448 219 25504
rect 275 25448 343 25504
rect 399 25448 467 25504
rect 523 25448 591 25504
rect 647 25448 715 25504
rect 771 25448 839 25504
rect 895 25448 1000 25504
rect 0 25380 1000 25448
rect 0 25324 95 25380
rect 151 25324 219 25380
rect 275 25324 343 25380
rect 399 25324 467 25380
rect 523 25324 591 25380
rect 647 25324 715 25380
rect 771 25324 839 25380
rect 895 25324 1000 25380
rect 0 25314 1000 25324
rect 0 25200 200 25314
rect 800 25200 1000 25314
rect 0 24894 200 25000
rect 800 24894 1000 25000
rect 0 24884 1000 24894
rect 0 24828 95 24884
rect 151 24828 219 24884
rect 275 24828 343 24884
rect 399 24828 467 24884
rect 523 24828 591 24884
rect 647 24828 715 24884
rect 771 24828 839 24884
rect 895 24828 1000 24884
rect 0 24760 1000 24828
rect 0 24704 95 24760
rect 151 24704 219 24760
rect 275 24704 343 24760
rect 399 24704 467 24760
rect 523 24704 591 24760
rect 647 24704 715 24760
rect 771 24704 839 24760
rect 895 24704 1000 24760
rect 0 24636 1000 24704
rect 0 24580 95 24636
rect 151 24580 219 24636
rect 275 24580 343 24636
rect 399 24580 467 24636
rect 523 24580 591 24636
rect 647 24580 715 24636
rect 771 24580 839 24636
rect 895 24580 1000 24636
rect 0 24512 1000 24580
rect 0 24456 95 24512
rect 151 24456 219 24512
rect 275 24456 343 24512
rect 399 24456 467 24512
rect 523 24456 591 24512
rect 647 24456 715 24512
rect 771 24456 839 24512
rect 895 24456 1000 24512
rect 0 24388 1000 24456
rect 0 24332 95 24388
rect 151 24332 219 24388
rect 275 24332 343 24388
rect 399 24332 467 24388
rect 523 24332 591 24388
rect 647 24332 715 24388
rect 771 24332 839 24388
rect 895 24332 1000 24388
rect 0 24264 1000 24332
rect 0 24208 95 24264
rect 151 24208 219 24264
rect 275 24208 343 24264
rect 399 24208 467 24264
rect 523 24208 591 24264
rect 647 24208 715 24264
rect 771 24208 839 24264
rect 895 24208 1000 24264
rect 0 24140 1000 24208
rect 0 24084 95 24140
rect 151 24084 219 24140
rect 275 24084 343 24140
rect 399 24084 467 24140
rect 523 24084 591 24140
rect 647 24084 715 24140
rect 771 24084 839 24140
rect 895 24084 1000 24140
rect 0 24016 1000 24084
rect 0 23960 95 24016
rect 151 23960 219 24016
rect 275 23960 343 24016
rect 399 23960 467 24016
rect 523 23960 591 24016
rect 647 23960 715 24016
rect 771 23960 839 24016
rect 895 23960 1000 24016
rect 0 23892 1000 23960
rect 0 23836 95 23892
rect 151 23836 219 23892
rect 275 23836 343 23892
rect 399 23836 467 23892
rect 523 23836 591 23892
rect 647 23836 715 23892
rect 771 23836 839 23892
rect 895 23836 1000 23892
rect 0 23768 1000 23836
rect 0 23712 95 23768
rect 151 23712 219 23768
rect 275 23712 343 23768
rect 399 23712 467 23768
rect 523 23712 591 23768
rect 647 23712 715 23768
rect 771 23712 839 23768
rect 895 23712 1000 23768
rect 0 23702 1000 23712
rect 0 23600 200 23702
rect 800 23600 1000 23702
rect 0 23307 200 23400
rect 800 23307 1000 23400
rect 0 23297 1000 23307
rect 0 23241 94 23297
rect 150 23241 218 23297
rect 274 23241 342 23297
rect 398 23241 466 23297
rect 522 23241 590 23297
rect 646 23241 714 23297
rect 770 23241 838 23297
rect 894 23241 1000 23297
rect 0 23173 1000 23241
rect 0 23117 94 23173
rect 150 23117 218 23173
rect 274 23117 342 23173
rect 398 23117 466 23173
rect 522 23117 590 23173
rect 646 23117 714 23173
rect 770 23117 838 23173
rect 894 23117 1000 23173
rect 0 23049 1000 23117
rect 0 22993 94 23049
rect 150 22993 218 23049
rect 274 22993 342 23049
rect 398 22993 466 23049
rect 522 22993 590 23049
rect 646 22993 714 23049
rect 770 22993 838 23049
rect 894 22993 1000 23049
rect 0 22925 1000 22993
rect 0 22869 94 22925
rect 150 22869 218 22925
rect 274 22869 342 22925
rect 398 22869 466 22925
rect 522 22869 590 22925
rect 646 22869 714 22925
rect 770 22869 838 22925
rect 894 22869 1000 22925
rect 0 22801 1000 22869
rect 0 22745 94 22801
rect 150 22745 218 22801
rect 274 22745 342 22801
rect 398 22745 466 22801
rect 522 22745 590 22801
rect 646 22745 714 22801
rect 770 22745 838 22801
rect 894 22745 1000 22801
rect 0 22677 1000 22745
rect 0 22621 94 22677
rect 150 22621 218 22677
rect 274 22621 342 22677
rect 398 22621 466 22677
rect 522 22621 590 22677
rect 646 22621 714 22677
rect 770 22621 838 22677
rect 894 22621 1000 22677
rect 0 22553 1000 22621
rect 0 22497 94 22553
rect 150 22497 218 22553
rect 274 22497 342 22553
rect 398 22497 466 22553
rect 522 22497 590 22553
rect 646 22497 714 22553
rect 770 22497 838 22553
rect 894 22497 1000 22553
rect 0 22429 1000 22497
rect 0 22373 94 22429
rect 150 22373 218 22429
rect 274 22373 342 22429
rect 398 22373 466 22429
rect 522 22373 590 22429
rect 646 22373 714 22429
rect 770 22373 838 22429
rect 894 22373 1000 22429
rect 0 22305 1000 22373
rect 0 22249 94 22305
rect 150 22249 218 22305
rect 274 22249 342 22305
rect 398 22249 466 22305
rect 522 22249 590 22305
rect 646 22249 714 22305
rect 770 22249 838 22305
rect 894 22249 1000 22305
rect 0 22181 1000 22249
rect 0 22125 94 22181
rect 150 22125 218 22181
rect 274 22125 342 22181
rect 398 22125 466 22181
rect 522 22125 590 22181
rect 646 22125 714 22181
rect 770 22125 838 22181
rect 894 22125 1000 22181
rect 0 22057 1000 22125
rect 0 22001 94 22057
rect 150 22001 218 22057
rect 274 22001 342 22057
rect 398 22001 466 22057
rect 522 22001 590 22057
rect 646 22001 714 22057
rect 770 22001 838 22057
rect 894 22001 1000 22057
rect 0 21933 1000 22001
rect 0 21877 94 21933
rect 150 21877 218 21933
rect 274 21877 342 21933
rect 398 21877 466 21933
rect 522 21877 590 21933
rect 646 21877 714 21933
rect 770 21877 838 21933
rect 894 21877 1000 21933
rect 0 21809 1000 21877
rect 0 21753 94 21809
rect 150 21753 218 21809
rect 274 21753 342 21809
rect 398 21753 466 21809
rect 522 21753 590 21809
rect 646 21753 714 21809
rect 770 21753 838 21809
rect 894 21753 1000 21809
rect 0 21685 1000 21753
rect 0 21629 94 21685
rect 150 21629 218 21685
rect 274 21629 342 21685
rect 398 21629 466 21685
rect 522 21629 590 21685
rect 646 21629 714 21685
rect 770 21629 838 21685
rect 894 21629 1000 21685
rect 0 21561 1000 21629
rect 0 21505 94 21561
rect 150 21505 218 21561
rect 274 21505 342 21561
rect 398 21505 466 21561
rect 522 21505 590 21561
rect 646 21505 714 21561
rect 770 21505 838 21561
rect 894 21505 1000 21561
rect 0 21437 1000 21505
rect 0 21381 94 21437
rect 150 21381 218 21437
rect 274 21381 342 21437
rect 398 21381 466 21437
rect 522 21381 590 21437
rect 646 21381 714 21437
rect 770 21381 838 21437
rect 894 21381 1000 21437
rect 0 21313 1000 21381
rect 0 21257 94 21313
rect 150 21257 218 21313
rect 274 21257 342 21313
rect 398 21257 466 21313
rect 522 21257 590 21313
rect 646 21257 714 21313
rect 770 21257 838 21313
rect 894 21257 1000 21313
rect 0 21189 1000 21257
rect 0 21133 94 21189
rect 150 21133 218 21189
rect 274 21133 342 21189
rect 398 21133 466 21189
rect 522 21133 590 21189
rect 646 21133 714 21189
rect 770 21133 838 21189
rect 894 21133 1000 21189
rect 0 21065 1000 21133
rect 0 21009 94 21065
rect 150 21009 218 21065
rect 274 21009 342 21065
rect 398 21009 466 21065
rect 522 21009 590 21065
rect 646 21009 714 21065
rect 770 21009 838 21065
rect 894 21009 1000 21065
rect 0 20941 1000 21009
rect 0 20885 94 20941
rect 150 20885 218 20941
rect 274 20885 342 20941
rect 398 20885 466 20941
rect 522 20885 590 20941
rect 646 20885 714 20941
rect 770 20885 838 20941
rect 894 20885 1000 20941
rect 0 20817 1000 20885
rect 0 20761 94 20817
rect 150 20761 218 20817
rect 274 20761 342 20817
rect 398 20761 466 20817
rect 522 20761 590 20817
rect 646 20761 714 20817
rect 770 20761 838 20817
rect 894 20761 1000 20817
rect 0 20693 1000 20761
rect 0 20637 94 20693
rect 150 20637 218 20693
rect 274 20637 342 20693
rect 398 20637 466 20693
rect 522 20637 590 20693
rect 646 20637 714 20693
rect 770 20637 838 20693
rect 894 20637 1000 20693
rect 0 20569 1000 20637
rect 0 20513 94 20569
rect 150 20513 218 20569
rect 274 20513 342 20569
rect 398 20513 466 20569
rect 522 20513 590 20569
rect 646 20513 714 20569
rect 770 20513 838 20569
rect 894 20513 1000 20569
rect 0 20503 1000 20513
rect 0 20400 200 20503
rect 800 20400 1000 20503
rect 0 20096 200 20200
rect 800 20096 1000 20200
rect 0 20086 1000 20096
rect 0 20030 94 20086
rect 150 20030 218 20086
rect 274 20030 342 20086
rect 398 20030 466 20086
rect 522 20030 590 20086
rect 646 20030 714 20086
rect 770 20030 838 20086
rect 894 20030 1000 20086
rect 0 19962 1000 20030
rect 0 19906 94 19962
rect 150 19906 218 19962
rect 274 19906 342 19962
rect 398 19906 466 19962
rect 522 19906 590 19962
rect 646 19906 714 19962
rect 770 19906 838 19962
rect 894 19906 1000 19962
rect 0 19838 1000 19906
rect 0 19782 94 19838
rect 150 19782 218 19838
rect 274 19782 342 19838
rect 398 19782 466 19838
rect 522 19782 590 19838
rect 646 19782 714 19838
rect 770 19782 838 19838
rect 894 19782 1000 19838
rect 0 19714 1000 19782
rect 0 19658 94 19714
rect 150 19658 218 19714
rect 274 19658 342 19714
rect 398 19658 466 19714
rect 522 19658 590 19714
rect 646 19658 714 19714
rect 770 19658 838 19714
rect 894 19658 1000 19714
rect 0 19590 1000 19658
rect 0 19534 94 19590
rect 150 19534 218 19590
rect 274 19534 342 19590
rect 398 19534 466 19590
rect 522 19534 590 19590
rect 646 19534 714 19590
rect 770 19534 838 19590
rect 894 19534 1000 19590
rect 0 19466 1000 19534
rect 0 19410 94 19466
rect 150 19410 218 19466
rect 274 19410 342 19466
rect 398 19410 466 19466
rect 522 19410 590 19466
rect 646 19410 714 19466
rect 770 19410 838 19466
rect 894 19410 1000 19466
rect 0 19342 1000 19410
rect 0 19286 94 19342
rect 150 19286 218 19342
rect 274 19286 342 19342
rect 398 19286 466 19342
rect 522 19286 590 19342
rect 646 19286 714 19342
rect 770 19286 838 19342
rect 894 19286 1000 19342
rect 0 19218 1000 19286
rect 0 19162 94 19218
rect 150 19162 218 19218
rect 274 19162 342 19218
rect 398 19162 466 19218
rect 522 19162 590 19218
rect 646 19162 714 19218
rect 770 19162 838 19218
rect 894 19162 1000 19218
rect 0 19094 1000 19162
rect 0 19038 94 19094
rect 150 19038 218 19094
rect 274 19038 342 19094
rect 398 19038 466 19094
rect 522 19038 590 19094
rect 646 19038 714 19094
rect 770 19038 838 19094
rect 894 19038 1000 19094
rect 0 18970 1000 19038
rect 0 18914 94 18970
rect 150 18914 218 18970
rect 274 18914 342 18970
rect 398 18914 466 18970
rect 522 18914 590 18970
rect 646 18914 714 18970
rect 770 18914 838 18970
rect 894 18914 1000 18970
rect 0 18846 1000 18914
rect 0 18790 94 18846
rect 150 18790 218 18846
rect 274 18790 342 18846
rect 398 18790 466 18846
rect 522 18790 590 18846
rect 646 18790 714 18846
rect 770 18790 838 18846
rect 894 18790 1000 18846
rect 0 18722 1000 18790
rect 0 18666 94 18722
rect 150 18666 218 18722
rect 274 18666 342 18722
rect 398 18666 466 18722
rect 522 18666 590 18722
rect 646 18666 714 18722
rect 770 18666 838 18722
rect 894 18666 1000 18722
rect 0 18598 1000 18666
rect 0 18542 94 18598
rect 150 18542 218 18598
rect 274 18542 342 18598
rect 398 18542 466 18598
rect 522 18542 590 18598
rect 646 18542 714 18598
rect 770 18542 838 18598
rect 894 18542 1000 18598
rect 0 18474 1000 18542
rect 0 18418 94 18474
rect 150 18418 218 18474
rect 274 18418 342 18474
rect 398 18418 466 18474
rect 522 18418 590 18474
rect 646 18418 714 18474
rect 770 18418 838 18474
rect 894 18418 1000 18474
rect 0 18350 1000 18418
rect 0 18294 94 18350
rect 150 18294 218 18350
rect 274 18294 342 18350
rect 398 18294 466 18350
rect 522 18294 590 18350
rect 646 18294 714 18350
rect 770 18294 838 18350
rect 894 18294 1000 18350
rect 0 18226 1000 18294
rect 0 18170 94 18226
rect 150 18170 218 18226
rect 274 18170 342 18226
rect 398 18170 466 18226
rect 522 18170 590 18226
rect 646 18170 714 18226
rect 770 18170 838 18226
rect 894 18170 1000 18226
rect 0 18102 1000 18170
rect 0 18046 94 18102
rect 150 18046 218 18102
rect 274 18046 342 18102
rect 398 18046 466 18102
rect 522 18046 590 18102
rect 646 18046 714 18102
rect 770 18046 838 18102
rect 894 18046 1000 18102
rect 0 17978 1000 18046
rect 0 17922 94 17978
rect 150 17922 218 17978
rect 274 17922 342 17978
rect 398 17922 466 17978
rect 522 17922 590 17978
rect 646 17922 714 17978
rect 770 17922 838 17978
rect 894 17922 1000 17978
rect 0 17854 1000 17922
rect 0 17798 94 17854
rect 150 17798 218 17854
rect 274 17798 342 17854
rect 398 17798 466 17854
rect 522 17798 590 17854
rect 646 17798 714 17854
rect 770 17798 838 17854
rect 894 17798 1000 17854
rect 0 17730 1000 17798
rect 0 17674 94 17730
rect 150 17674 218 17730
rect 274 17674 342 17730
rect 398 17674 466 17730
rect 522 17674 590 17730
rect 646 17674 714 17730
rect 770 17674 838 17730
rect 894 17674 1000 17730
rect 0 17606 1000 17674
rect 0 17550 94 17606
rect 150 17550 218 17606
rect 274 17550 342 17606
rect 398 17550 466 17606
rect 522 17550 590 17606
rect 646 17550 714 17606
rect 770 17550 838 17606
rect 894 17550 1000 17606
rect 0 17482 1000 17550
rect 0 17426 94 17482
rect 150 17426 218 17482
rect 274 17426 342 17482
rect 398 17426 466 17482
rect 522 17426 590 17482
rect 646 17426 714 17482
rect 770 17426 838 17482
rect 894 17426 1000 17482
rect 0 17358 1000 17426
rect 0 17302 94 17358
rect 150 17302 218 17358
rect 274 17302 342 17358
rect 398 17302 466 17358
rect 522 17302 590 17358
rect 646 17302 714 17358
rect 770 17302 838 17358
rect 894 17302 1000 17358
rect 0 17292 1000 17302
rect 0 17200 200 17292
rect 800 17200 1000 17292
rect 0 16923 200 17000
rect 800 16923 1000 17000
rect 0 16913 1000 16923
rect 0 16857 94 16913
rect 150 16857 218 16913
rect 274 16857 342 16913
rect 398 16857 466 16913
rect 522 16857 590 16913
rect 646 16857 714 16913
rect 770 16857 838 16913
rect 894 16857 1000 16913
rect 0 16789 1000 16857
rect 0 16733 94 16789
rect 150 16733 218 16789
rect 274 16733 342 16789
rect 398 16733 466 16789
rect 522 16733 590 16789
rect 646 16733 714 16789
rect 770 16733 838 16789
rect 894 16733 1000 16789
rect 0 16665 1000 16733
rect 0 16609 94 16665
rect 150 16609 218 16665
rect 274 16609 342 16665
rect 398 16609 466 16665
rect 522 16609 590 16665
rect 646 16609 714 16665
rect 770 16609 838 16665
rect 894 16609 1000 16665
rect 0 16541 1000 16609
rect 0 16485 94 16541
rect 150 16485 218 16541
rect 274 16485 342 16541
rect 398 16485 466 16541
rect 522 16485 590 16541
rect 646 16485 714 16541
rect 770 16485 838 16541
rect 894 16485 1000 16541
rect 0 16417 1000 16485
rect 0 16361 94 16417
rect 150 16361 218 16417
rect 274 16361 342 16417
rect 398 16361 466 16417
rect 522 16361 590 16417
rect 646 16361 714 16417
rect 770 16361 838 16417
rect 894 16361 1000 16417
rect 0 16293 1000 16361
rect 0 16237 94 16293
rect 150 16237 218 16293
rect 274 16237 342 16293
rect 398 16237 466 16293
rect 522 16237 590 16293
rect 646 16237 714 16293
rect 770 16237 838 16293
rect 894 16237 1000 16293
rect 0 16169 1000 16237
rect 0 16113 94 16169
rect 150 16113 218 16169
rect 274 16113 342 16169
rect 398 16113 466 16169
rect 522 16113 590 16169
rect 646 16113 714 16169
rect 770 16113 838 16169
rect 894 16113 1000 16169
rect 0 16045 1000 16113
rect 0 15989 94 16045
rect 150 15989 218 16045
rect 274 15989 342 16045
rect 398 15989 466 16045
rect 522 15989 590 16045
rect 646 15989 714 16045
rect 770 15989 838 16045
rect 894 15989 1000 16045
rect 0 15921 1000 15989
rect 0 15865 94 15921
rect 150 15865 218 15921
rect 274 15865 342 15921
rect 398 15865 466 15921
rect 522 15865 590 15921
rect 646 15865 714 15921
rect 770 15865 838 15921
rect 894 15865 1000 15921
rect 0 15797 1000 15865
rect 0 15741 94 15797
rect 150 15741 218 15797
rect 274 15741 342 15797
rect 398 15741 466 15797
rect 522 15741 590 15797
rect 646 15741 714 15797
rect 770 15741 838 15797
rect 894 15741 1000 15797
rect 0 15673 1000 15741
rect 0 15617 94 15673
rect 150 15617 218 15673
rect 274 15617 342 15673
rect 398 15617 466 15673
rect 522 15617 590 15673
rect 646 15617 714 15673
rect 770 15617 838 15673
rect 894 15617 1000 15673
rect 0 15549 1000 15617
rect 0 15493 94 15549
rect 150 15493 218 15549
rect 274 15493 342 15549
rect 398 15493 466 15549
rect 522 15493 590 15549
rect 646 15493 714 15549
rect 770 15493 838 15549
rect 894 15493 1000 15549
rect 0 15425 1000 15493
rect 0 15369 94 15425
rect 150 15369 218 15425
rect 274 15369 342 15425
rect 398 15369 466 15425
rect 522 15369 590 15425
rect 646 15369 714 15425
rect 770 15369 838 15425
rect 894 15369 1000 15425
rect 0 15301 1000 15369
rect 0 15245 94 15301
rect 150 15245 218 15301
rect 274 15245 342 15301
rect 398 15245 466 15301
rect 522 15245 590 15301
rect 646 15245 714 15301
rect 770 15245 838 15301
rect 894 15245 1000 15301
rect 0 15177 1000 15245
rect 0 15121 94 15177
rect 150 15121 218 15177
rect 274 15121 342 15177
rect 398 15121 466 15177
rect 522 15121 590 15177
rect 646 15121 714 15177
rect 770 15121 838 15177
rect 894 15121 1000 15177
rect 0 15053 1000 15121
rect 0 14997 94 15053
rect 150 14997 218 15053
rect 274 14997 342 15053
rect 398 14997 466 15053
rect 522 14997 590 15053
rect 646 14997 714 15053
rect 770 14997 838 15053
rect 894 14997 1000 15053
rect 0 14929 1000 14997
rect 0 14873 94 14929
rect 150 14873 218 14929
rect 274 14873 342 14929
rect 398 14873 466 14929
rect 522 14873 590 14929
rect 646 14873 714 14929
rect 770 14873 838 14929
rect 894 14873 1000 14929
rect 0 14805 1000 14873
rect 0 14749 94 14805
rect 150 14749 218 14805
rect 274 14749 342 14805
rect 398 14749 466 14805
rect 522 14749 590 14805
rect 646 14749 714 14805
rect 770 14749 838 14805
rect 894 14749 1000 14805
rect 0 14681 1000 14749
rect 0 14625 94 14681
rect 150 14625 218 14681
rect 274 14625 342 14681
rect 398 14625 466 14681
rect 522 14625 590 14681
rect 646 14625 714 14681
rect 770 14625 838 14681
rect 894 14625 1000 14681
rect 0 14557 1000 14625
rect 0 14501 94 14557
rect 150 14501 218 14557
rect 274 14501 342 14557
rect 398 14501 466 14557
rect 522 14501 590 14557
rect 646 14501 714 14557
rect 770 14501 838 14557
rect 894 14501 1000 14557
rect 0 14433 1000 14501
rect 0 14377 94 14433
rect 150 14377 218 14433
rect 274 14377 342 14433
rect 398 14377 466 14433
rect 522 14377 590 14433
rect 646 14377 714 14433
rect 770 14377 838 14433
rect 894 14377 1000 14433
rect 0 14309 1000 14377
rect 0 14253 94 14309
rect 150 14253 218 14309
rect 274 14253 342 14309
rect 398 14253 466 14309
rect 522 14253 590 14309
rect 646 14253 714 14309
rect 770 14253 838 14309
rect 894 14253 1000 14309
rect 0 14185 1000 14253
rect 0 14129 94 14185
rect 150 14129 218 14185
rect 274 14129 342 14185
rect 398 14129 466 14185
rect 522 14129 590 14185
rect 646 14129 714 14185
rect 770 14129 838 14185
rect 894 14129 1000 14185
rect 0 14119 1000 14129
rect 0 14000 200 14119
rect 800 14000 1000 14119
<< via3 >>
rect 94 69573 150 69629
rect 218 69573 274 69629
rect 342 69573 398 69629
rect 466 69573 522 69629
rect 590 69573 646 69629
rect 714 69573 770 69629
rect 838 69573 894 69629
rect 94 69449 150 69505
rect 218 69449 274 69505
rect 342 69449 398 69505
rect 466 69449 522 69505
rect 590 69449 646 69505
rect 714 69449 770 69505
rect 838 69449 894 69505
rect 94 69325 150 69381
rect 218 69325 274 69381
rect 342 69325 398 69381
rect 466 69325 522 69381
rect 590 69325 646 69381
rect 714 69325 770 69381
rect 838 69325 894 69381
rect 94 69201 150 69257
rect 218 69201 274 69257
rect 342 69201 398 69257
rect 466 69201 522 69257
rect 590 69201 646 69257
rect 714 69201 770 69257
rect 838 69201 894 69257
rect 94 69077 150 69133
rect 218 69077 274 69133
rect 342 69077 398 69133
rect 466 69077 522 69133
rect 590 69077 646 69133
rect 714 69077 770 69133
rect 838 69077 894 69133
rect 94 68953 150 69009
rect 218 68953 274 69009
rect 342 68953 398 69009
rect 466 68953 522 69009
rect 590 68953 646 69009
rect 714 68953 770 69009
rect 838 68953 894 69009
rect 94 68829 150 68885
rect 218 68829 274 68885
rect 342 68829 398 68885
rect 466 68829 522 68885
rect 590 68829 646 68885
rect 714 68829 770 68885
rect 838 68829 894 68885
rect 94 68705 150 68761
rect 218 68705 274 68761
rect 342 68705 398 68761
rect 466 68705 522 68761
rect 590 68705 646 68761
rect 714 68705 770 68761
rect 838 68705 894 68761
rect 94 68581 150 68637
rect 218 68581 274 68637
rect 342 68581 398 68637
rect 466 68581 522 68637
rect 590 68581 646 68637
rect 714 68581 770 68637
rect 838 68581 894 68637
rect 94 68457 150 68513
rect 218 68457 274 68513
rect 342 68457 398 68513
rect 466 68457 522 68513
rect 590 68457 646 68513
rect 714 68457 770 68513
rect 838 68457 894 68513
rect 94 68028 150 68084
rect 218 68028 274 68084
rect 342 68028 398 68084
rect 466 68028 522 68084
rect 590 68028 646 68084
rect 714 68028 770 68084
rect 838 68028 894 68084
rect 94 67904 150 67960
rect 218 67904 274 67960
rect 342 67904 398 67960
rect 466 67904 522 67960
rect 590 67904 646 67960
rect 714 67904 770 67960
rect 838 67904 894 67960
rect 94 67780 150 67836
rect 218 67780 274 67836
rect 342 67780 398 67836
rect 466 67780 522 67836
rect 590 67780 646 67836
rect 714 67780 770 67836
rect 838 67780 894 67836
rect 94 67656 150 67712
rect 218 67656 274 67712
rect 342 67656 398 67712
rect 466 67656 522 67712
rect 590 67656 646 67712
rect 714 67656 770 67712
rect 838 67656 894 67712
rect 94 67532 150 67588
rect 218 67532 274 67588
rect 342 67532 398 67588
rect 466 67532 522 67588
rect 590 67532 646 67588
rect 714 67532 770 67588
rect 838 67532 894 67588
rect 94 67408 150 67464
rect 218 67408 274 67464
rect 342 67408 398 67464
rect 466 67408 522 67464
rect 590 67408 646 67464
rect 714 67408 770 67464
rect 838 67408 894 67464
rect 94 67284 150 67340
rect 218 67284 274 67340
rect 342 67284 398 67340
rect 466 67284 522 67340
rect 590 67284 646 67340
rect 714 67284 770 67340
rect 838 67284 894 67340
rect 94 67160 150 67216
rect 218 67160 274 67216
rect 342 67160 398 67216
rect 466 67160 522 67216
rect 590 67160 646 67216
rect 714 67160 770 67216
rect 838 67160 894 67216
rect 94 67036 150 67092
rect 218 67036 274 67092
rect 342 67036 398 67092
rect 466 67036 522 67092
rect 590 67036 646 67092
rect 714 67036 770 67092
rect 838 67036 894 67092
rect 94 66912 150 66968
rect 218 66912 274 66968
rect 342 66912 398 66968
rect 466 66912 522 66968
rect 590 66912 646 66968
rect 714 66912 770 66968
rect 838 66912 894 66968
rect 94 66421 150 66477
rect 218 66421 274 66477
rect 342 66421 398 66477
rect 466 66421 522 66477
rect 590 66421 646 66477
rect 714 66421 770 66477
rect 838 66421 894 66477
rect 94 66297 150 66353
rect 218 66297 274 66353
rect 342 66297 398 66353
rect 466 66297 522 66353
rect 590 66297 646 66353
rect 714 66297 770 66353
rect 838 66297 894 66353
rect 94 66173 150 66229
rect 218 66173 274 66229
rect 342 66173 398 66229
rect 466 66173 522 66229
rect 590 66173 646 66229
rect 714 66173 770 66229
rect 838 66173 894 66229
rect 94 66049 150 66105
rect 218 66049 274 66105
rect 342 66049 398 66105
rect 466 66049 522 66105
rect 590 66049 646 66105
rect 714 66049 770 66105
rect 838 66049 894 66105
rect 94 65925 150 65981
rect 218 65925 274 65981
rect 342 65925 398 65981
rect 466 65925 522 65981
rect 590 65925 646 65981
rect 714 65925 770 65981
rect 838 65925 894 65981
rect 94 65801 150 65857
rect 218 65801 274 65857
rect 342 65801 398 65857
rect 466 65801 522 65857
rect 590 65801 646 65857
rect 714 65801 770 65857
rect 838 65801 894 65857
rect 94 65677 150 65733
rect 218 65677 274 65733
rect 342 65677 398 65733
rect 466 65677 522 65733
rect 590 65677 646 65733
rect 714 65677 770 65733
rect 838 65677 894 65733
rect 94 65553 150 65609
rect 218 65553 274 65609
rect 342 65553 398 65609
rect 466 65553 522 65609
rect 590 65553 646 65609
rect 714 65553 770 65609
rect 838 65553 894 65609
rect 94 65429 150 65485
rect 218 65429 274 65485
rect 342 65429 398 65485
rect 466 65429 522 65485
rect 590 65429 646 65485
rect 714 65429 770 65485
rect 838 65429 894 65485
rect 94 65305 150 65361
rect 218 65305 274 65361
rect 342 65305 398 65361
rect 466 65305 522 65361
rect 590 65305 646 65361
rect 714 65305 770 65361
rect 838 65305 894 65361
rect 94 64830 150 64886
rect 218 64830 274 64886
rect 342 64830 398 64886
rect 466 64830 522 64886
rect 590 64830 646 64886
rect 714 64830 770 64886
rect 838 64830 894 64886
rect 94 64706 150 64762
rect 218 64706 274 64762
rect 342 64706 398 64762
rect 466 64706 522 64762
rect 590 64706 646 64762
rect 714 64706 770 64762
rect 838 64706 894 64762
rect 94 64582 150 64638
rect 218 64582 274 64638
rect 342 64582 398 64638
rect 466 64582 522 64638
rect 590 64582 646 64638
rect 714 64582 770 64638
rect 838 64582 894 64638
rect 94 64458 150 64514
rect 218 64458 274 64514
rect 342 64458 398 64514
rect 466 64458 522 64514
rect 590 64458 646 64514
rect 714 64458 770 64514
rect 838 64458 894 64514
rect 94 64334 150 64390
rect 218 64334 274 64390
rect 342 64334 398 64390
rect 466 64334 522 64390
rect 590 64334 646 64390
rect 714 64334 770 64390
rect 838 64334 894 64390
rect 94 64210 150 64266
rect 218 64210 274 64266
rect 342 64210 398 64266
rect 466 64210 522 64266
rect 590 64210 646 64266
rect 714 64210 770 64266
rect 838 64210 894 64266
rect 94 64086 150 64142
rect 218 64086 274 64142
rect 342 64086 398 64142
rect 466 64086 522 64142
rect 590 64086 646 64142
rect 714 64086 770 64142
rect 838 64086 894 64142
rect 94 63962 150 64018
rect 218 63962 274 64018
rect 342 63962 398 64018
rect 466 63962 522 64018
rect 590 63962 646 64018
rect 714 63962 770 64018
rect 838 63962 894 64018
rect 94 63838 150 63894
rect 218 63838 274 63894
rect 342 63838 398 63894
rect 466 63838 522 63894
rect 590 63838 646 63894
rect 714 63838 770 63894
rect 838 63838 894 63894
rect 94 63714 150 63770
rect 218 63714 274 63770
rect 342 63714 398 63770
rect 466 63714 522 63770
rect 590 63714 646 63770
rect 714 63714 770 63770
rect 838 63714 894 63770
rect 94 63224 150 63280
rect 218 63224 274 63280
rect 342 63224 398 63280
rect 466 63224 522 63280
rect 590 63224 646 63280
rect 714 63224 770 63280
rect 838 63224 894 63280
rect 94 63100 150 63156
rect 218 63100 274 63156
rect 342 63100 398 63156
rect 466 63100 522 63156
rect 590 63100 646 63156
rect 714 63100 770 63156
rect 838 63100 894 63156
rect 94 62976 150 63032
rect 218 62976 274 63032
rect 342 62976 398 63032
rect 466 62976 522 63032
rect 590 62976 646 63032
rect 714 62976 770 63032
rect 838 62976 894 63032
rect 94 62852 150 62908
rect 218 62852 274 62908
rect 342 62852 398 62908
rect 466 62852 522 62908
rect 590 62852 646 62908
rect 714 62852 770 62908
rect 838 62852 894 62908
rect 94 62728 150 62784
rect 218 62728 274 62784
rect 342 62728 398 62784
rect 466 62728 522 62784
rect 590 62728 646 62784
rect 714 62728 770 62784
rect 838 62728 894 62784
rect 94 62604 150 62660
rect 218 62604 274 62660
rect 342 62604 398 62660
rect 466 62604 522 62660
rect 590 62604 646 62660
rect 714 62604 770 62660
rect 838 62604 894 62660
rect 94 62480 150 62536
rect 218 62480 274 62536
rect 342 62480 398 62536
rect 466 62480 522 62536
rect 590 62480 646 62536
rect 714 62480 770 62536
rect 838 62480 894 62536
rect 94 62356 150 62412
rect 218 62356 274 62412
rect 342 62356 398 62412
rect 466 62356 522 62412
rect 590 62356 646 62412
rect 714 62356 770 62412
rect 838 62356 894 62412
rect 94 62232 150 62288
rect 218 62232 274 62288
rect 342 62232 398 62288
rect 466 62232 522 62288
rect 590 62232 646 62288
rect 714 62232 770 62288
rect 838 62232 894 62288
rect 94 62108 150 62164
rect 218 62108 274 62164
rect 342 62108 398 62164
rect 466 62108 522 62164
rect 590 62108 646 62164
rect 714 62108 770 62164
rect 838 62108 894 62164
rect 94 61638 150 61694
rect 218 61638 274 61694
rect 342 61638 398 61694
rect 466 61638 522 61694
rect 590 61638 646 61694
rect 714 61638 770 61694
rect 838 61638 894 61694
rect 94 61514 150 61570
rect 218 61514 274 61570
rect 342 61514 398 61570
rect 466 61514 522 61570
rect 590 61514 646 61570
rect 714 61514 770 61570
rect 838 61514 894 61570
rect 94 61390 150 61446
rect 218 61390 274 61446
rect 342 61390 398 61446
rect 466 61390 522 61446
rect 590 61390 646 61446
rect 714 61390 770 61446
rect 838 61390 894 61446
rect 94 61266 150 61322
rect 218 61266 274 61322
rect 342 61266 398 61322
rect 466 61266 522 61322
rect 590 61266 646 61322
rect 714 61266 770 61322
rect 838 61266 894 61322
rect 94 61142 150 61198
rect 218 61142 274 61198
rect 342 61142 398 61198
rect 466 61142 522 61198
rect 590 61142 646 61198
rect 714 61142 770 61198
rect 838 61142 894 61198
rect 94 61018 150 61074
rect 218 61018 274 61074
rect 342 61018 398 61074
rect 466 61018 522 61074
rect 590 61018 646 61074
rect 714 61018 770 61074
rect 838 61018 894 61074
rect 94 60894 150 60950
rect 218 60894 274 60950
rect 342 60894 398 60950
rect 466 60894 522 60950
rect 590 60894 646 60950
rect 714 60894 770 60950
rect 838 60894 894 60950
rect 94 60770 150 60826
rect 218 60770 274 60826
rect 342 60770 398 60826
rect 466 60770 522 60826
rect 590 60770 646 60826
rect 714 60770 770 60826
rect 838 60770 894 60826
rect 94 60646 150 60702
rect 218 60646 274 60702
rect 342 60646 398 60702
rect 466 60646 522 60702
rect 590 60646 646 60702
rect 714 60646 770 60702
rect 838 60646 894 60702
rect 94 60522 150 60578
rect 218 60522 274 60578
rect 342 60522 398 60578
rect 466 60522 522 60578
rect 590 60522 646 60578
rect 714 60522 770 60578
rect 838 60522 894 60578
rect 94 60046 150 60102
rect 218 60046 274 60102
rect 342 60046 398 60102
rect 466 60046 522 60102
rect 590 60046 646 60102
rect 714 60046 770 60102
rect 838 60046 894 60102
rect 94 59922 150 59978
rect 218 59922 274 59978
rect 342 59922 398 59978
rect 466 59922 522 59978
rect 590 59922 646 59978
rect 714 59922 770 59978
rect 838 59922 894 59978
rect 94 59798 150 59854
rect 218 59798 274 59854
rect 342 59798 398 59854
rect 466 59798 522 59854
rect 590 59798 646 59854
rect 714 59798 770 59854
rect 838 59798 894 59854
rect 94 59674 150 59730
rect 218 59674 274 59730
rect 342 59674 398 59730
rect 466 59674 522 59730
rect 590 59674 646 59730
rect 714 59674 770 59730
rect 838 59674 894 59730
rect 94 59550 150 59606
rect 218 59550 274 59606
rect 342 59550 398 59606
rect 466 59550 522 59606
rect 590 59550 646 59606
rect 714 59550 770 59606
rect 838 59550 894 59606
rect 94 59426 150 59482
rect 218 59426 274 59482
rect 342 59426 398 59482
rect 466 59426 522 59482
rect 590 59426 646 59482
rect 714 59426 770 59482
rect 838 59426 894 59482
rect 94 59302 150 59358
rect 218 59302 274 59358
rect 342 59302 398 59358
rect 466 59302 522 59358
rect 590 59302 646 59358
rect 714 59302 770 59358
rect 838 59302 894 59358
rect 94 59178 150 59234
rect 218 59178 274 59234
rect 342 59178 398 59234
rect 466 59178 522 59234
rect 590 59178 646 59234
rect 714 59178 770 59234
rect 838 59178 894 59234
rect 94 59054 150 59110
rect 218 59054 274 59110
rect 342 59054 398 59110
rect 466 59054 522 59110
rect 590 59054 646 59110
rect 714 59054 770 59110
rect 838 59054 894 59110
rect 94 58930 150 58986
rect 218 58930 274 58986
rect 342 58930 398 58986
rect 466 58930 522 58986
rect 590 58930 646 58986
rect 714 58930 770 58986
rect 838 58930 894 58986
rect 94 58429 150 58485
rect 218 58429 274 58485
rect 342 58429 398 58485
rect 466 58429 522 58485
rect 590 58429 646 58485
rect 714 58429 770 58485
rect 838 58429 894 58485
rect 94 58305 150 58361
rect 218 58305 274 58361
rect 342 58305 398 58361
rect 466 58305 522 58361
rect 590 58305 646 58361
rect 714 58305 770 58361
rect 838 58305 894 58361
rect 94 58181 150 58237
rect 218 58181 274 58237
rect 342 58181 398 58237
rect 466 58181 522 58237
rect 590 58181 646 58237
rect 714 58181 770 58237
rect 838 58181 894 58237
rect 94 58057 150 58113
rect 218 58057 274 58113
rect 342 58057 398 58113
rect 466 58057 522 58113
rect 590 58057 646 58113
rect 714 58057 770 58113
rect 838 58057 894 58113
rect 94 57933 150 57989
rect 218 57933 274 57989
rect 342 57933 398 57989
rect 466 57933 522 57989
rect 590 57933 646 57989
rect 714 57933 770 57989
rect 838 57933 894 57989
rect 94 57809 150 57865
rect 218 57809 274 57865
rect 342 57809 398 57865
rect 466 57809 522 57865
rect 590 57809 646 57865
rect 714 57809 770 57865
rect 838 57809 894 57865
rect 94 57685 150 57741
rect 218 57685 274 57741
rect 342 57685 398 57741
rect 466 57685 522 57741
rect 590 57685 646 57741
rect 714 57685 770 57741
rect 838 57685 894 57741
rect 94 57561 150 57617
rect 218 57561 274 57617
rect 342 57561 398 57617
rect 466 57561 522 57617
rect 590 57561 646 57617
rect 714 57561 770 57617
rect 838 57561 894 57617
rect 94 57437 150 57493
rect 218 57437 274 57493
rect 342 57437 398 57493
rect 466 57437 522 57493
rect 590 57437 646 57493
rect 714 57437 770 57493
rect 838 57437 894 57493
rect 94 57313 150 57369
rect 218 57313 274 57369
rect 342 57313 398 57369
rect 466 57313 522 57369
rect 590 57313 646 57369
rect 714 57313 770 57369
rect 838 57313 894 57369
rect 94 56836 150 56892
rect 218 56836 274 56892
rect 342 56836 398 56892
rect 466 56836 522 56892
rect 590 56836 646 56892
rect 714 56836 770 56892
rect 838 56836 894 56892
rect 94 56712 150 56768
rect 218 56712 274 56768
rect 342 56712 398 56768
rect 466 56712 522 56768
rect 590 56712 646 56768
rect 714 56712 770 56768
rect 838 56712 894 56768
rect 94 56588 150 56644
rect 218 56588 274 56644
rect 342 56588 398 56644
rect 466 56588 522 56644
rect 590 56588 646 56644
rect 714 56588 770 56644
rect 838 56588 894 56644
rect 94 56464 150 56520
rect 218 56464 274 56520
rect 342 56464 398 56520
rect 466 56464 522 56520
rect 590 56464 646 56520
rect 714 56464 770 56520
rect 838 56464 894 56520
rect 94 56340 150 56396
rect 218 56340 274 56396
rect 342 56340 398 56396
rect 466 56340 522 56396
rect 590 56340 646 56396
rect 714 56340 770 56396
rect 838 56340 894 56396
rect 94 56216 150 56272
rect 218 56216 274 56272
rect 342 56216 398 56272
rect 466 56216 522 56272
rect 590 56216 646 56272
rect 714 56216 770 56272
rect 838 56216 894 56272
rect 94 56092 150 56148
rect 218 56092 274 56148
rect 342 56092 398 56148
rect 466 56092 522 56148
rect 590 56092 646 56148
rect 714 56092 770 56148
rect 838 56092 894 56148
rect 94 55968 150 56024
rect 218 55968 274 56024
rect 342 55968 398 56024
rect 466 55968 522 56024
rect 590 55968 646 56024
rect 714 55968 770 56024
rect 838 55968 894 56024
rect 94 55844 150 55900
rect 218 55844 274 55900
rect 342 55844 398 55900
rect 466 55844 522 55900
rect 590 55844 646 55900
rect 714 55844 770 55900
rect 838 55844 894 55900
rect 94 55720 150 55776
rect 218 55720 274 55776
rect 342 55720 398 55776
rect 466 55720 522 55776
rect 590 55720 646 55776
rect 714 55720 770 55776
rect 838 55720 894 55776
rect 94 55232 150 55288
rect 218 55232 274 55288
rect 342 55232 398 55288
rect 466 55232 522 55288
rect 590 55232 646 55288
rect 714 55232 770 55288
rect 838 55232 894 55288
rect 94 55108 150 55164
rect 218 55108 274 55164
rect 342 55108 398 55164
rect 466 55108 522 55164
rect 590 55108 646 55164
rect 714 55108 770 55164
rect 838 55108 894 55164
rect 94 54984 150 55040
rect 218 54984 274 55040
rect 342 54984 398 55040
rect 466 54984 522 55040
rect 590 54984 646 55040
rect 714 54984 770 55040
rect 838 54984 894 55040
rect 94 54860 150 54916
rect 218 54860 274 54916
rect 342 54860 398 54916
rect 466 54860 522 54916
rect 590 54860 646 54916
rect 714 54860 770 54916
rect 838 54860 894 54916
rect 94 54736 150 54792
rect 218 54736 274 54792
rect 342 54736 398 54792
rect 466 54736 522 54792
rect 590 54736 646 54792
rect 714 54736 770 54792
rect 838 54736 894 54792
rect 94 54612 150 54668
rect 218 54612 274 54668
rect 342 54612 398 54668
rect 466 54612 522 54668
rect 590 54612 646 54668
rect 714 54612 770 54668
rect 838 54612 894 54668
rect 94 54488 150 54544
rect 218 54488 274 54544
rect 342 54488 398 54544
rect 466 54488 522 54544
rect 590 54488 646 54544
rect 714 54488 770 54544
rect 838 54488 894 54544
rect 94 54364 150 54420
rect 218 54364 274 54420
rect 342 54364 398 54420
rect 466 54364 522 54420
rect 590 54364 646 54420
rect 714 54364 770 54420
rect 838 54364 894 54420
rect 94 54240 150 54296
rect 218 54240 274 54296
rect 342 54240 398 54296
rect 466 54240 522 54296
rect 590 54240 646 54296
rect 714 54240 770 54296
rect 838 54240 894 54296
rect 94 54116 150 54172
rect 218 54116 274 54172
rect 342 54116 398 54172
rect 466 54116 522 54172
rect 590 54116 646 54172
rect 714 54116 770 54172
rect 838 54116 894 54172
rect 94 53626 150 53682
rect 218 53626 274 53682
rect 342 53626 398 53682
rect 466 53626 522 53682
rect 590 53626 646 53682
rect 714 53626 770 53682
rect 838 53626 894 53682
rect 94 53502 150 53558
rect 218 53502 274 53558
rect 342 53502 398 53558
rect 466 53502 522 53558
rect 590 53502 646 53558
rect 714 53502 770 53558
rect 838 53502 894 53558
rect 94 53378 150 53434
rect 218 53378 274 53434
rect 342 53378 398 53434
rect 466 53378 522 53434
rect 590 53378 646 53434
rect 714 53378 770 53434
rect 838 53378 894 53434
rect 94 53254 150 53310
rect 218 53254 274 53310
rect 342 53254 398 53310
rect 466 53254 522 53310
rect 590 53254 646 53310
rect 714 53254 770 53310
rect 838 53254 894 53310
rect 94 53130 150 53186
rect 218 53130 274 53186
rect 342 53130 398 53186
rect 466 53130 522 53186
rect 590 53130 646 53186
rect 714 53130 770 53186
rect 838 53130 894 53186
rect 94 53006 150 53062
rect 218 53006 274 53062
rect 342 53006 398 53062
rect 466 53006 522 53062
rect 590 53006 646 53062
rect 714 53006 770 53062
rect 838 53006 894 53062
rect 94 52882 150 52938
rect 218 52882 274 52938
rect 342 52882 398 52938
rect 466 52882 522 52938
rect 590 52882 646 52938
rect 714 52882 770 52938
rect 838 52882 894 52938
rect 94 52758 150 52814
rect 218 52758 274 52814
rect 342 52758 398 52814
rect 466 52758 522 52814
rect 590 52758 646 52814
rect 714 52758 770 52814
rect 838 52758 894 52814
rect 94 52634 150 52690
rect 218 52634 274 52690
rect 342 52634 398 52690
rect 466 52634 522 52690
rect 590 52634 646 52690
rect 714 52634 770 52690
rect 838 52634 894 52690
rect 94 52510 150 52566
rect 218 52510 274 52566
rect 342 52510 398 52566
rect 466 52510 522 52566
rect 590 52510 646 52566
rect 714 52510 770 52566
rect 838 52510 894 52566
rect 94 52023 150 52079
rect 218 52023 274 52079
rect 342 52023 398 52079
rect 466 52023 522 52079
rect 590 52023 646 52079
rect 714 52023 770 52079
rect 838 52023 894 52079
rect 94 51899 150 51955
rect 218 51899 274 51955
rect 342 51899 398 51955
rect 466 51899 522 51955
rect 590 51899 646 51955
rect 714 51899 770 51955
rect 838 51899 894 51955
rect 94 51775 150 51831
rect 218 51775 274 51831
rect 342 51775 398 51831
rect 466 51775 522 51831
rect 590 51775 646 51831
rect 714 51775 770 51831
rect 838 51775 894 51831
rect 94 51651 150 51707
rect 218 51651 274 51707
rect 342 51651 398 51707
rect 466 51651 522 51707
rect 590 51651 646 51707
rect 714 51651 770 51707
rect 838 51651 894 51707
rect 94 51527 150 51583
rect 218 51527 274 51583
rect 342 51527 398 51583
rect 466 51527 522 51583
rect 590 51527 646 51583
rect 714 51527 770 51583
rect 838 51527 894 51583
rect 94 51403 150 51459
rect 218 51403 274 51459
rect 342 51403 398 51459
rect 466 51403 522 51459
rect 590 51403 646 51459
rect 714 51403 770 51459
rect 838 51403 894 51459
rect 94 51279 150 51335
rect 218 51279 274 51335
rect 342 51279 398 51335
rect 466 51279 522 51335
rect 590 51279 646 51335
rect 714 51279 770 51335
rect 838 51279 894 51335
rect 94 51155 150 51211
rect 218 51155 274 51211
rect 342 51155 398 51211
rect 466 51155 522 51211
rect 590 51155 646 51211
rect 714 51155 770 51211
rect 838 51155 894 51211
rect 94 51031 150 51087
rect 218 51031 274 51087
rect 342 51031 398 51087
rect 466 51031 522 51087
rect 590 51031 646 51087
rect 714 51031 770 51087
rect 838 51031 894 51087
rect 94 50907 150 50963
rect 218 50907 274 50963
rect 342 50907 398 50963
rect 466 50907 522 50963
rect 590 50907 646 50963
rect 714 50907 770 50963
rect 838 50907 894 50963
rect 95 50424 151 50480
rect 219 50424 275 50480
rect 343 50424 399 50480
rect 467 50424 523 50480
rect 591 50424 647 50480
rect 715 50424 771 50480
rect 839 50424 895 50480
rect 95 50300 151 50356
rect 219 50300 275 50356
rect 343 50300 399 50356
rect 467 50300 523 50356
rect 591 50300 647 50356
rect 715 50300 771 50356
rect 839 50300 895 50356
rect 95 50176 151 50232
rect 219 50176 275 50232
rect 343 50176 399 50232
rect 467 50176 523 50232
rect 591 50176 647 50232
rect 715 50176 771 50232
rect 839 50176 895 50232
rect 95 50052 151 50108
rect 219 50052 275 50108
rect 343 50052 399 50108
rect 467 50052 523 50108
rect 591 50052 647 50108
rect 715 50052 771 50108
rect 839 50052 895 50108
rect 95 49928 151 49984
rect 219 49928 275 49984
rect 343 49928 399 49984
rect 467 49928 523 49984
rect 591 49928 647 49984
rect 715 49928 771 49984
rect 839 49928 895 49984
rect 95 49804 151 49860
rect 219 49804 275 49860
rect 343 49804 399 49860
rect 467 49804 523 49860
rect 591 49804 647 49860
rect 715 49804 771 49860
rect 839 49804 895 49860
rect 95 49680 151 49736
rect 219 49680 275 49736
rect 343 49680 399 49736
rect 467 49680 523 49736
rect 591 49680 647 49736
rect 715 49680 771 49736
rect 839 49680 895 49736
rect 95 49556 151 49612
rect 219 49556 275 49612
rect 343 49556 399 49612
rect 467 49556 523 49612
rect 591 49556 647 49612
rect 715 49556 771 49612
rect 839 49556 895 49612
rect 95 49432 151 49488
rect 219 49432 275 49488
rect 343 49432 399 49488
rect 467 49432 523 49488
rect 591 49432 647 49488
rect 715 49432 771 49488
rect 839 49432 895 49488
rect 95 49308 151 49364
rect 219 49308 275 49364
rect 343 49308 399 49364
rect 467 49308 523 49364
rect 591 49308 647 49364
rect 715 49308 771 49364
rect 839 49308 895 49364
rect 94 48837 150 48893
rect 218 48837 274 48893
rect 342 48837 398 48893
rect 466 48837 522 48893
rect 590 48837 646 48893
rect 714 48837 770 48893
rect 838 48837 894 48893
rect 94 48713 150 48769
rect 218 48713 274 48769
rect 342 48713 398 48769
rect 466 48713 522 48769
rect 590 48713 646 48769
rect 714 48713 770 48769
rect 838 48713 894 48769
rect 94 48589 150 48645
rect 218 48589 274 48645
rect 342 48589 398 48645
rect 466 48589 522 48645
rect 590 48589 646 48645
rect 714 48589 770 48645
rect 838 48589 894 48645
rect 94 48465 150 48521
rect 218 48465 274 48521
rect 342 48465 398 48521
rect 466 48465 522 48521
rect 590 48465 646 48521
rect 714 48465 770 48521
rect 838 48465 894 48521
rect 94 48341 150 48397
rect 218 48341 274 48397
rect 342 48341 398 48397
rect 466 48341 522 48397
rect 590 48341 646 48397
rect 714 48341 770 48397
rect 838 48341 894 48397
rect 94 48217 150 48273
rect 218 48217 274 48273
rect 342 48217 398 48273
rect 466 48217 522 48273
rect 590 48217 646 48273
rect 714 48217 770 48273
rect 838 48217 894 48273
rect 94 48093 150 48149
rect 218 48093 274 48149
rect 342 48093 398 48149
rect 466 48093 522 48149
rect 590 48093 646 48149
rect 714 48093 770 48149
rect 838 48093 894 48149
rect 94 47969 150 48025
rect 218 47969 274 48025
rect 342 47969 398 48025
rect 466 47969 522 48025
rect 590 47969 646 48025
rect 714 47969 770 48025
rect 838 47969 894 48025
rect 94 47845 150 47901
rect 218 47845 274 47901
rect 342 47845 398 47901
rect 466 47845 522 47901
rect 590 47845 646 47901
rect 714 47845 770 47901
rect 838 47845 894 47901
rect 94 47721 150 47777
rect 218 47721 274 47777
rect 342 47721 398 47777
rect 466 47721 522 47777
rect 590 47721 646 47777
rect 714 47721 770 47777
rect 838 47721 894 47777
rect 94 47597 150 47653
rect 218 47597 274 47653
rect 342 47597 398 47653
rect 466 47597 522 47653
rect 590 47597 646 47653
rect 714 47597 770 47653
rect 838 47597 894 47653
rect 94 47473 150 47529
rect 218 47473 274 47529
rect 342 47473 398 47529
rect 466 47473 522 47529
rect 590 47473 646 47529
rect 714 47473 770 47529
rect 838 47473 894 47529
rect 94 47349 150 47405
rect 218 47349 274 47405
rect 342 47349 398 47405
rect 466 47349 522 47405
rect 590 47349 646 47405
rect 714 47349 770 47405
rect 838 47349 894 47405
rect 94 47225 150 47281
rect 218 47225 274 47281
rect 342 47225 398 47281
rect 466 47225 522 47281
rect 590 47225 646 47281
rect 714 47225 770 47281
rect 838 47225 894 47281
rect 94 47101 150 47157
rect 218 47101 274 47157
rect 342 47101 398 47157
rect 466 47101 522 47157
rect 590 47101 646 47157
rect 714 47101 770 47157
rect 838 47101 894 47157
rect 94 46977 150 47033
rect 218 46977 274 47033
rect 342 46977 398 47033
rect 466 46977 522 47033
rect 590 46977 646 47033
rect 714 46977 770 47033
rect 838 46977 894 47033
rect 94 46853 150 46909
rect 218 46853 274 46909
rect 342 46853 398 46909
rect 466 46853 522 46909
rect 590 46853 646 46909
rect 714 46853 770 46909
rect 838 46853 894 46909
rect 94 46729 150 46785
rect 218 46729 274 46785
rect 342 46729 398 46785
rect 466 46729 522 46785
rect 590 46729 646 46785
rect 714 46729 770 46785
rect 838 46729 894 46785
rect 94 46605 150 46661
rect 218 46605 274 46661
rect 342 46605 398 46661
rect 466 46605 522 46661
rect 590 46605 646 46661
rect 714 46605 770 46661
rect 838 46605 894 46661
rect 94 46481 150 46537
rect 218 46481 274 46537
rect 342 46481 398 46537
rect 466 46481 522 46537
rect 590 46481 646 46537
rect 714 46481 770 46537
rect 838 46481 894 46537
rect 94 46357 150 46413
rect 218 46357 274 46413
rect 342 46357 398 46413
rect 466 46357 522 46413
rect 590 46357 646 46413
rect 714 46357 770 46413
rect 838 46357 894 46413
rect 94 46233 150 46289
rect 218 46233 274 46289
rect 342 46233 398 46289
rect 466 46233 522 46289
rect 590 46233 646 46289
rect 714 46233 770 46289
rect 838 46233 894 46289
rect 94 46109 150 46165
rect 218 46109 274 46165
rect 342 46109 398 46165
rect 466 46109 522 46165
rect 590 46109 646 46165
rect 714 46109 770 46165
rect 838 46109 894 46165
rect 94 45641 150 45697
rect 218 45641 274 45697
rect 342 45641 398 45697
rect 466 45641 522 45697
rect 590 45641 646 45697
rect 714 45641 770 45697
rect 838 45641 894 45697
rect 94 45517 150 45573
rect 218 45517 274 45573
rect 342 45517 398 45573
rect 466 45517 522 45573
rect 590 45517 646 45573
rect 714 45517 770 45573
rect 838 45517 894 45573
rect 94 45393 150 45449
rect 218 45393 274 45449
rect 342 45393 398 45449
rect 466 45393 522 45449
rect 590 45393 646 45449
rect 714 45393 770 45449
rect 838 45393 894 45449
rect 94 45269 150 45325
rect 218 45269 274 45325
rect 342 45269 398 45325
rect 466 45269 522 45325
rect 590 45269 646 45325
rect 714 45269 770 45325
rect 838 45269 894 45325
rect 94 45145 150 45201
rect 218 45145 274 45201
rect 342 45145 398 45201
rect 466 45145 522 45201
rect 590 45145 646 45201
rect 714 45145 770 45201
rect 838 45145 894 45201
rect 94 45021 150 45077
rect 218 45021 274 45077
rect 342 45021 398 45077
rect 466 45021 522 45077
rect 590 45021 646 45077
rect 714 45021 770 45077
rect 838 45021 894 45077
rect 94 44897 150 44953
rect 218 44897 274 44953
rect 342 44897 398 44953
rect 466 44897 522 44953
rect 590 44897 646 44953
rect 714 44897 770 44953
rect 838 44897 894 44953
rect 94 44773 150 44829
rect 218 44773 274 44829
rect 342 44773 398 44829
rect 466 44773 522 44829
rect 590 44773 646 44829
rect 714 44773 770 44829
rect 838 44773 894 44829
rect 94 44649 150 44705
rect 218 44649 274 44705
rect 342 44649 398 44705
rect 466 44649 522 44705
rect 590 44649 646 44705
rect 714 44649 770 44705
rect 838 44649 894 44705
rect 94 44525 150 44581
rect 218 44525 274 44581
rect 342 44525 398 44581
rect 466 44525 522 44581
rect 590 44525 646 44581
rect 714 44525 770 44581
rect 838 44525 894 44581
rect 94 44401 150 44457
rect 218 44401 274 44457
rect 342 44401 398 44457
rect 466 44401 522 44457
rect 590 44401 646 44457
rect 714 44401 770 44457
rect 838 44401 894 44457
rect 94 44277 150 44333
rect 218 44277 274 44333
rect 342 44277 398 44333
rect 466 44277 522 44333
rect 590 44277 646 44333
rect 714 44277 770 44333
rect 838 44277 894 44333
rect 94 44153 150 44209
rect 218 44153 274 44209
rect 342 44153 398 44209
rect 466 44153 522 44209
rect 590 44153 646 44209
rect 714 44153 770 44209
rect 838 44153 894 44209
rect 94 44029 150 44085
rect 218 44029 274 44085
rect 342 44029 398 44085
rect 466 44029 522 44085
rect 590 44029 646 44085
rect 714 44029 770 44085
rect 838 44029 894 44085
rect 94 43905 150 43961
rect 218 43905 274 43961
rect 342 43905 398 43961
rect 466 43905 522 43961
rect 590 43905 646 43961
rect 714 43905 770 43961
rect 838 43905 894 43961
rect 94 43781 150 43837
rect 218 43781 274 43837
rect 342 43781 398 43837
rect 466 43781 522 43837
rect 590 43781 646 43837
rect 714 43781 770 43837
rect 838 43781 894 43837
rect 94 43657 150 43713
rect 218 43657 274 43713
rect 342 43657 398 43713
rect 466 43657 522 43713
rect 590 43657 646 43713
rect 714 43657 770 43713
rect 838 43657 894 43713
rect 94 43533 150 43589
rect 218 43533 274 43589
rect 342 43533 398 43589
rect 466 43533 522 43589
rect 590 43533 646 43589
rect 714 43533 770 43589
rect 838 43533 894 43589
rect 94 43409 150 43465
rect 218 43409 274 43465
rect 342 43409 398 43465
rect 466 43409 522 43465
rect 590 43409 646 43465
rect 714 43409 770 43465
rect 838 43409 894 43465
rect 94 43285 150 43341
rect 218 43285 274 43341
rect 342 43285 398 43341
rect 466 43285 522 43341
rect 590 43285 646 43341
rect 714 43285 770 43341
rect 838 43285 894 43341
rect 94 43161 150 43217
rect 218 43161 274 43217
rect 342 43161 398 43217
rect 466 43161 522 43217
rect 590 43161 646 43217
rect 714 43161 770 43217
rect 838 43161 894 43217
rect 94 43037 150 43093
rect 218 43037 274 43093
rect 342 43037 398 43093
rect 466 43037 522 43093
rect 590 43037 646 43093
rect 714 43037 770 43093
rect 838 43037 894 43093
rect 94 42913 150 42969
rect 218 42913 274 42969
rect 342 42913 398 42969
rect 466 42913 522 42969
rect 590 42913 646 42969
rect 714 42913 770 42969
rect 838 42913 894 42969
rect 95 42428 151 42484
rect 219 42428 275 42484
rect 343 42428 399 42484
rect 467 42428 523 42484
rect 591 42428 647 42484
rect 715 42428 771 42484
rect 839 42428 895 42484
rect 95 42304 151 42360
rect 219 42304 275 42360
rect 343 42304 399 42360
rect 467 42304 523 42360
rect 591 42304 647 42360
rect 715 42304 771 42360
rect 839 42304 895 42360
rect 95 42180 151 42236
rect 219 42180 275 42236
rect 343 42180 399 42236
rect 467 42180 523 42236
rect 591 42180 647 42236
rect 715 42180 771 42236
rect 839 42180 895 42236
rect 95 42056 151 42112
rect 219 42056 275 42112
rect 343 42056 399 42112
rect 467 42056 523 42112
rect 591 42056 647 42112
rect 715 42056 771 42112
rect 839 42056 895 42112
rect 95 41932 151 41988
rect 219 41932 275 41988
rect 343 41932 399 41988
rect 467 41932 523 41988
rect 591 41932 647 41988
rect 715 41932 771 41988
rect 839 41932 895 41988
rect 95 41808 151 41864
rect 219 41808 275 41864
rect 343 41808 399 41864
rect 467 41808 523 41864
rect 591 41808 647 41864
rect 715 41808 771 41864
rect 839 41808 895 41864
rect 95 41684 151 41740
rect 219 41684 275 41740
rect 343 41684 399 41740
rect 467 41684 523 41740
rect 591 41684 647 41740
rect 715 41684 771 41740
rect 839 41684 895 41740
rect 95 41560 151 41616
rect 219 41560 275 41616
rect 343 41560 399 41616
rect 467 41560 523 41616
rect 591 41560 647 41616
rect 715 41560 771 41616
rect 839 41560 895 41616
rect 95 41436 151 41492
rect 219 41436 275 41492
rect 343 41436 399 41492
rect 467 41436 523 41492
rect 591 41436 647 41492
rect 715 41436 771 41492
rect 839 41436 895 41492
rect 95 41312 151 41368
rect 219 41312 275 41368
rect 343 41312 399 41368
rect 467 41312 523 41368
rect 591 41312 647 41368
rect 715 41312 771 41368
rect 839 41312 895 41368
rect 95 40840 151 40896
rect 219 40840 275 40896
rect 343 40840 399 40896
rect 467 40840 523 40896
rect 591 40840 647 40896
rect 715 40840 771 40896
rect 839 40840 895 40896
rect 95 40716 151 40772
rect 219 40716 275 40772
rect 343 40716 399 40772
rect 467 40716 523 40772
rect 591 40716 647 40772
rect 715 40716 771 40772
rect 839 40716 895 40772
rect 95 40592 151 40648
rect 219 40592 275 40648
rect 343 40592 399 40648
rect 467 40592 523 40648
rect 591 40592 647 40648
rect 715 40592 771 40648
rect 839 40592 895 40648
rect 95 40468 151 40524
rect 219 40468 275 40524
rect 343 40468 399 40524
rect 467 40468 523 40524
rect 591 40468 647 40524
rect 715 40468 771 40524
rect 839 40468 895 40524
rect 95 40344 151 40400
rect 219 40344 275 40400
rect 343 40344 399 40400
rect 467 40344 523 40400
rect 591 40344 647 40400
rect 715 40344 771 40400
rect 839 40344 895 40400
rect 95 40220 151 40276
rect 219 40220 275 40276
rect 343 40220 399 40276
rect 467 40220 523 40276
rect 591 40220 647 40276
rect 715 40220 771 40276
rect 839 40220 895 40276
rect 95 40096 151 40152
rect 219 40096 275 40152
rect 343 40096 399 40152
rect 467 40096 523 40152
rect 591 40096 647 40152
rect 715 40096 771 40152
rect 839 40096 895 40152
rect 95 39972 151 40028
rect 219 39972 275 40028
rect 343 39972 399 40028
rect 467 39972 523 40028
rect 591 39972 647 40028
rect 715 39972 771 40028
rect 839 39972 895 40028
rect 95 39848 151 39904
rect 219 39848 275 39904
rect 343 39848 399 39904
rect 467 39848 523 39904
rect 591 39848 647 39904
rect 715 39848 771 39904
rect 839 39848 895 39904
rect 95 39724 151 39780
rect 219 39724 275 39780
rect 343 39724 399 39780
rect 467 39724 523 39780
rect 591 39724 647 39780
rect 715 39724 771 39780
rect 839 39724 895 39780
rect 94 39248 150 39304
rect 218 39248 274 39304
rect 342 39248 398 39304
rect 466 39248 522 39304
rect 590 39248 646 39304
rect 714 39248 770 39304
rect 838 39248 894 39304
rect 94 39124 150 39180
rect 218 39124 274 39180
rect 342 39124 398 39180
rect 466 39124 522 39180
rect 590 39124 646 39180
rect 714 39124 770 39180
rect 838 39124 894 39180
rect 94 39000 150 39056
rect 218 39000 274 39056
rect 342 39000 398 39056
rect 466 39000 522 39056
rect 590 39000 646 39056
rect 714 39000 770 39056
rect 838 39000 894 39056
rect 94 38876 150 38932
rect 218 38876 274 38932
rect 342 38876 398 38932
rect 466 38876 522 38932
rect 590 38876 646 38932
rect 714 38876 770 38932
rect 838 38876 894 38932
rect 94 38752 150 38808
rect 218 38752 274 38808
rect 342 38752 398 38808
rect 466 38752 522 38808
rect 590 38752 646 38808
rect 714 38752 770 38808
rect 838 38752 894 38808
rect 94 38628 150 38684
rect 218 38628 274 38684
rect 342 38628 398 38684
rect 466 38628 522 38684
rect 590 38628 646 38684
rect 714 38628 770 38684
rect 838 38628 894 38684
rect 94 38504 150 38560
rect 218 38504 274 38560
rect 342 38504 398 38560
rect 466 38504 522 38560
rect 590 38504 646 38560
rect 714 38504 770 38560
rect 838 38504 894 38560
rect 94 38380 150 38436
rect 218 38380 274 38436
rect 342 38380 398 38436
rect 466 38380 522 38436
rect 590 38380 646 38436
rect 714 38380 770 38436
rect 838 38380 894 38436
rect 94 38256 150 38312
rect 218 38256 274 38312
rect 342 38256 398 38312
rect 466 38256 522 38312
rect 590 38256 646 38312
rect 714 38256 770 38312
rect 838 38256 894 38312
rect 94 38132 150 38188
rect 218 38132 274 38188
rect 342 38132 398 38188
rect 466 38132 522 38188
rect 590 38132 646 38188
rect 714 38132 770 38188
rect 838 38132 894 38188
rect 94 38008 150 38064
rect 218 38008 274 38064
rect 342 38008 398 38064
rect 466 38008 522 38064
rect 590 38008 646 38064
rect 714 38008 770 38064
rect 838 38008 894 38064
rect 94 37884 150 37940
rect 218 37884 274 37940
rect 342 37884 398 37940
rect 466 37884 522 37940
rect 590 37884 646 37940
rect 714 37884 770 37940
rect 838 37884 894 37940
rect 94 37760 150 37816
rect 218 37760 274 37816
rect 342 37760 398 37816
rect 466 37760 522 37816
rect 590 37760 646 37816
rect 714 37760 770 37816
rect 838 37760 894 37816
rect 94 37636 150 37692
rect 218 37636 274 37692
rect 342 37636 398 37692
rect 466 37636 522 37692
rect 590 37636 646 37692
rect 714 37636 770 37692
rect 838 37636 894 37692
rect 94 37512 150 37568
rect 218 37512 274 37568
rect 342 37512 398 37568
rect 466 37512 522 37568
rect 590 37512 646 37568
rect 714 37512 770 37568
rect 838 37512 894 37568
rect 94 37388 150 37444
rect 218 37388 274 37444
rect 342 37388 398 37444
rect 466 37388 522 37444
rect 590 37388 646 37444
rect 714 37388 770 37444
rect 838 37388 894 37444
rect 94 37264 150 37320
rect 218 37264 274 37320
rect 342 37264 398 37320
rect 466 37264 522 37320
rect 590 37264 646 37320
rect 714 37264 770 37320
rect 838 37264 894 37320
rect 94 37140 150 37196
rect 218 37140 274 37196
rect 342 37140 398 37196
rect 466 37140 522 37196
rect 590 37140 646 37196
rect 714 37140 770 37196
rect 838 37140 894 37196
rect 94 37016 150 37072
rect 218 37016 274 37072
rect 342 37016 398 37072
rect 466 37016 522 37072
rect 590 37016 646 37072
rect 714 37016 770 37072
rect 838 37016 894 37072
rect 94 36892 150 36948
rect 218 36892 274 36948
rect 342 36892 398 36948
rect 466 36892 522 36948
rect 590 36892 646 36948
rect 714 36892 770 36948
rect 838 36892 894 36948
rect 94 36768 150 36824
rect 218 36768 274 36824
rect 342 36768 398 36824
rect 466 36768 522 36824
rect 590 36768 646 36824
rect 714 36768 770 36824
rect 838 36768 894 36824
rect 94 36644 150 36700
rect 218 36644 274 36700
rect 342 36644 398 36700
rect 466 36644 522 36700
rect 590 36644 646 36700
rect 714 36644 770 36700
rect 838 36644 894 36700
rect 94 36520 150 36576
rect 218 36520 274 36576
rect 342 36520 398 36576
rect 466 36520 522 36576
rect 590 36520 646 36576
rect 714 36520 770 36576
rect 838 36520 894 36576
rect 94 36038 150 36094
rect 218 36038 274 36094
rect 342 36038 398 36094
rect 466 36038 522 36094
rect 590 36038 646 36094
rect 714 36038 770 36094
rect 838 36038 894 36094
rect 94 35914 150 35970
rect 218 35914 274 35970
rect 342 35914 398 35970
rect 466 35914 522 35970
rect 590 35914 646 35970
rect 714 35914 770 35970
rect 838 35914 894 35970
rect 94 35790 150 35846
rect 218 35790 274 35846
rect 342 35790 398 35846
rect 466 35790 522 35846
rect 590 35790 646 35846
rect 714 35790 770 35846
rect 838 35790 894 35846
rect 94 35666 150 35722
rect 218 35666 274 35722
rect 342 35666 398 35722
rect 466 35666 522 35722
rect 590 35666 646 35722
rect 714 35666 770 35722
rect 838 35666 894 35722
rect 94 35542 150 35598
rect 218 35542 274 35598
rect 342 35542 398 35598
rect 466 35542 522 35598
rect 590 35542 646 35598
rect 714 35542 770 35598
rect 838 35542 894 35598
rect 94 35418 150 35474
rect 218 35418 274 35474
rect 342 35418 398 35474
rect 466 35418 522 35474
rect 590 35418 646 35474
rect 714 35418 770 35474
rect 838 35418 894 35474
rect 94 35294 150 35350
rect 218 35294 274 35350
rect 342 35294 398 35350
rect 466 35294 522 35350
rect 590 35294 646 35350
rect 714 35294 770 35350
rect 838 35294 894 35350
rect 94 35170 150 35226
rect 218 35170 274 35226
rect 342 35170 398 35226
rect 466 35170 522 35226
rect 590 35170 646 35226
rect 714 35170 770 35226
rect 838 35170 894 35226
rect 94 35046 150 35102
rect 218 35046 274 35102
rect 342 35046 398 35102
rect 466 35046 522 35102
rect 590 35046 646 35102
rect 714 35046 770 35102
rect 838 35046 894 35102
rect 94 34922 150 34978
rect 218 34922 274 34978
rect 342 34922 398 34978
rect 466 34922 522 34978
rect 590 34922 646 34978
rect 714 34922 770 34978
rect 838 34922 894 34978
rect 94 34798 150 34854
rect 218 34798 274 34854
rect 342 34798 398 34854
rect 466 34798 522 34854
rect 590 34798 646 34854
rect 714 34798 770 34854
rect 838 34798 894 34854
rect 94 34674 150 34730
rect 218 34674 274 34730
rect 342 34674 398 34730
rect 466 34674 522 34730
rect 590 34674 646 34730
rect 714 34674 770 34730
rect 838 34674 894 34730
rect 94 34550 150 34606
rect 218 34550 274 34606
rect 342 34550 398 34606
rect 466 34550 522 34606
rect 590 34550 646 34606
rect 714 34550 770 34606
rect 838 34550 894 34606
rect 94 34426 150 34482
rect 218 34426 274 34482
rect 342 34426 398 34482
rect 466 34426 522 34482
rect 590 34426 646 34482
rect 714 34426 770 34482
rect 838 34426 894 34482
rect 94 34302 150 34358
rect 218 34302 274 34358
rect 342 34302 398 34358
rect 466 34302 522 34358
rect 590 34302 646 34358
rect 714 34302 770 34358
rect 838 34302 894 34358
rect 94 34178 150 34234
rect 218 34178 274 34234
rect 342 34178 398 34234
rect 466 34178 522 34234
rect 590 34178 646 34234
rect 714 34178 770 34234
rect 838 34178 894 34234
rect 94 34054 150 34110
rect 218 34054 274 34110
rect 342 34054 398 34110
rect 466 34054 522 34110
rect 590 34054 646 34110
rect 714 34054 770 34110
rect 838 34054 894 34110
rect 94 33930 150 33986
rect 218 33930 274 33986
rect 342 33930 398 33986
rect 466 33930 522 33986
rect 590 33930 646 33986
rect 714 33930 770 33986
rect 838 33930 894 33986
rect 94 33806 150 33862
rect 218 33806 274 33862
rect 342 33806 398 33862
rect 466 33806 522 33862
rect 590 33806 646 33862
rect 714 33806 770 33862
rect 838 33806 894 33862
rect 94 33682 150 33738
rect 218 33682 274 33738
rect 342 33682 398 33738
rect 466 33682 522 33738
rect 590 33682 646 33738
rect 714 33682 770 33738
rect 838 33682 894 33738
rect 94 33558 150 33614
rect 218 33558 274 33614
rect 342 33558 398 33614
rect 466 33558 522 33614
rect 590 33558 646 33614
rect 714 33558 770 33614
rect 838 33558 894 33614
rect 94 33434 150 33490
rect 218 33434 274 33490
rect 342 33434 398 33490
rect 466 33434 522 33490
rect 590 33434 646 33490
rect 714 33434 770 33490
rect 838 33434 894 33490
rect 94 33310 150 33366
rect 218 33310 274 33366
rect 342 33310 398 33366
rect 466 33310 522 33366
rect 590 33310 646 33366
rect 714 33310 770 33366
rect 838 33310 894 33366
rect 94 32846 150 32902
rect 218 32846 274 32902
rect 342 32846 398 32902
rect 466 32846 522 32902
rect 590 32846 646 32902
rect 714 32846 770 32902
rect 838 32846 894 32902
rect 94 32722 150 32778
rect 218 32722 274 32778
rect 342 32722 398 32778
rect 466 32722 522 32778
rect 590 32722 646 32778
rect 714 32722 770 32778
rect 838 32722 894 32778
rect 94 32598 150 32654
rect 218 32598 274 32654
rect 342 32598 398 32654
rect 466 32598 522 32654
rect 590 32598 646 32654
rect 714 32598 770 32654
rect 838 32598 894 32654
rect 94 32474 150 32530
rect 218 32474 274 32530
rect 342 32474 398 32530
rect 466 32474 522 32530
rect 590 32474 646 32530
rect 714 32474 770 32530
rect 838 32474 894 32530
rect 94 32350 150 32406
rect 218 32350 274 32406
rect 342 32350 398 32406
rect 466 32350 522 32406
rect 590 32350 646 32406
rect 714 32350 770 32406
rect 838 32350 894 32406
rect 94 32226 150 32282
rect 218 32226 274 32282
rect 342 32226 398 32282
rect 466 32226 522 32282
rect 590 32226 646 32282
rect 714 32226 770 32282
rect 838 32226 894 32282
rect 94 32102 150 32158
rect 218 32102 274 32158
rect 342 32102 398 32158
rect 466 32102 522 32158
rect 590 32102 646 32158
rect 714 32102 770 32158
rect 838 32102 894 32158
rect 94 31978 150 32034
rect 218 31978 274 32034
rect 342 31978 398 32034
rect 466 31978 522 32034
rect 590 31978 646 32034
rect 714 31978 770 32034
rect 838 31978 894 32034
rect 94 31854 150 31910
rect 218 31854 274 31910
rect 342 31854 398 31910
rect 466 31854 522 31910
rect 590 31854 646 31910
rect 714 31854 770 31910
rect 838 31854 894 31910
rect 94 31730 150 31786
rect 218 31730 274 31786
rect 342 31730 398 31786
rect 466 31730 522 31786
rect 590 31730 646 31786
rect 714 31730 770 31786
rect 838 31730 894 31786
rect 94 31606 150 31662
rect 218 31606 274 31662
rect 342 31606 398 31662
rect 466 31606 522 31662
rect 590 31606 646 31662
rect 714 31606 770 31662
rect 838 31606 894 31662
rect 94 31482 150 31538
rect 218 31482 274 31538
rect 342 31482 398 31538
rect 466 31482 522 31538
rect 590 31482 646 31538
rect 714 31482 770 31538
rect 838 31482 894 31538
rect 94 31358 150 31414
rect 218 31358 274 31414
rect 342 31358 398 31414
rect 466 31358 522 31414
rect 590 31358 646 31414
rect 714 31358 770 31414
rect 838 31358 894 31414
rect 94 31234 150 31290
rect 218 31234 274 31290
rect 342 31234 398 31290
rect 466 31234 522 31290
rect 590 31234 646 31290
rect 714 31234 770 31290
rect 838 31234 894 31290
rect 94 31110 150 31166
rect 218 31110 274 31166
rect 342 31110 398 31166
rect 466 31110 522 31166
rect 590 31110 646 31166
rect 714 31110 770 31166
rect 838 31110 894 31166
rect 94 30986 150 31042
rect 218 30986 274 31042
rect 342 30986 398 31042
rect 466 30986 522 31042
rect 590 30986 646 31042
rect 714 30986 770 31042
rect 838 30986 894 31042
rect 94 30862 150 30918
rect 218 30862 274 30918
rect 342 30862 398 30918
rect 466 30862 522 30918
rect 590 30862 646 30918
rect 714 30862 770 30918
rect 838 30862 894 30918
rect 94 30738 150 30794
rect 218 30738 274 30794
rect 342 30738 398 30794
rect 466 30738 522 30794
rect 590 30738 646 30794
rect 714 30738 770 30794
rect 838 30738 894 30794
rect 94 30614 150 30670
rect 218 30614 274 30670
rect 342 30614 398 30670
rect 466 30614 522 30670
rect 590 30614 646 30670
rect 714 30614 770 30670
rect 838 30614 894 30670
rect 94 30490 150 30546
rect 218 30490 274 30546
rect 342 30490 398 30546
rect 466 30490 522 30546
rect 590 30490 646 30546
rect 714 30490 770 30546
rect 838 30490 894 30546
rect 94 30366 150 30422
rect 218 30366 274 30422
rect 342 30366 398 30422
rect 466 30366 522 30422
rect 590 30366 646 30422
rect 714 30366 770 30422
rect 838 30366 894 30422
rect 94 30242 150 30298
rect 218 30242 274 30298
rect 342 30242 398 30298
rect 466 30242 522 30298
rect 590 30242 646 30298
rect 714 30242 770 30298
rect 838 30242 894 30298
rect 94 30118 150 30174
rect 218 30118 274 30174
rect 342 30118 398 30174
rect 466 30118 522 30174
rect 590 30118 646 30174
rect 714 30118 770 30174
rect 838 30118 894 30174
rect 94 29629 150 29685
rect 218 29629 274 29685
rect 342 29629 398 29685
rect 466 29629 522 29685
rect 590 29629 646 29685
rect 714 29629 770 29685
rect 838 29629 894 29685
rect 94 29505 150 29561
rect 218 29505 274 29561
rect 342 29505 398 29561
rect 466 29505 522 29561
rect 590 29505 646 29561
rect 714 29505 770 29561
rect 838 29505 894 29561
rect 94 29381 150 29437
rect 218 29381 274 29437
rect 342 29381 398 29437
rect 466 29381 522 29437
rect 590 29381 646 29437
rect 714 29381 770 29437
rect 838 29381 894 29437
rect 94 29257 150 29313
rect 218 29257 274 29313
rect 342 29257 398 29313
rect 466 29257 522 29313
rect 590 29257 646 29313
rect 714 29257 770 29313
rect 838 29257 894 29313
rect 94 29133 150 29189
rect 218 29133 274 29189
rect 342 29133 398 29189
rect 466 29133 522 29189
rect 590 29133 646 29189
rect 714 29133 770 29189
rect 838 29133 894 29189
rect 94 29009 150 29065
rect 218 29009 274 29065
rect 342 29009 398 29065
rect 466 29009 522 29065
rect 590 29009 646 29065
rect 714 29009 770 29065
rect 838 29009 894 29065
rect 94 28885 150 28941
rect 218 28885 274 28941
rect 342 28885 398 28941
rect 466 28885 522 28941
rect 590 28885 646 28941
rect 714 28885 770 28941
rect 838 28885 894 28941
rect 94 28761 150 28817
rect 218 28761 274 28817
rect 342 28761 398 28817
rect 466 28761 522 28817
rect 590 28761 646 28817
rect 714 28761 770 28817
rect 838 28761 894 28817
rect 94 28637 150 28693
rect 218 28637 274 28693
rect 342 28637 398 28693
rect 466 28637 522 28693
rect 590 28637 646 28693
rect 714 28637 770 28693
rect 838 28637 894 28693
rect 94 28513 150 28569
rect 218 28513 274 28569
rect 342 28513 398 28569
rect 466 28513 522 28569
rect 590 28513 646 28569
rect 714 28513 770 28569
rect 838 28513 894 28569
rect 94 28389 150 28445
rect 218 28389 274 28445
rect 342 28389 398 28445
rect 466 28389 522 28445
rect 590 28389 646 28445
rect 714 28389 770 28445
rect 838 28389 894 28445
rect 94 28265 150 28321
rect 218 28265 274 28321
rect 342 28265 398 28321
rect 466 28265 522 28321
rect 590 28265 646 28321
rect 714 28265 770 28321
rect 838 28265 894 28321
rect 94 28141 150 28197
rect 218 28141 274 28197
rect 342 28141 398 28197
rect 466 28141 522 28197
rect 590 28141 646 28197
rect 714 28141 770 28197
rect 838 28141 894 28197
rect 94 28017 150 28073
rect 218 28017 274 28073
rect 342 28017 398 28073
rect 466 28017 522 28073
rect 590 28017 646 28073
rect 714 28017 770 28073
rect 838 28017 894 28073
rect 94 27893 150 27949
rect 218 27893 274 27949
rect 342 27893 398 27949
rect 466 27893 522 27949
rect 590 27893 646 27949
rect 714 27893 770 27949
rect 838 27893 894 27949
rect 94 27769 150 27825
rect 218 27769 274 27825
rect 342 27769 398 27825
rect 466 27769 522 27825
rect 590 27769 646 27825
rect 714 27769 770 27825
rect 838 27769 894 27825
rect 94 27645 150 27701
rect 218 27645 274 27701
rect 342 27645 398 27701
rect 466 27645 522 27701
rect 590 27645 646 27701
rect 714 27645 770 27701
rect 838 27645 894 27701
rect 94 27521 150 27577
rect 218 27521 274 27577
rect 342 27521 398 27577
rect 466 27521 522 27577
rect 590 27521 646 27577
rect 714 27521 770 27577
rect 838 27521 894 27577
rect 94 27397 150 27453
rect 218 27397 274 27453
rect 342 27397 398 27453
rect 466 27397 522 27453
rect 590 27397 646 27453
rect 714 27397 770 27453
rect 838 27397 894 27453
rect 94 27273 150 27329
rect 218 27273 274 27329
rect 342 27273 398 27329
rect 466 27273 522 27329
rect 590 27273 646 27329
rect 714 27273 770 27329
rect 838 27273 894 27329
rect 94 27149 150 27205
rect 218 27149 274 27205
rect 342 27149 398 27205
rect 466 27149 522 27205
rect 590 27149 646 27205
rect 714 27149 770 27205
rect 838 27149 894 27205
rect 94 27025 150 27081
rect 218 27025 274 27081
rect 342 27025 398 27081
rect 466 27025 522 27081
rect 590 27025 646 27081
rect 714 27025 770 27081
rect 838 27025 894 27081
rect 94 26901 150 26957
rect 218 26901 274 26957
rect 342 26901 398 26957
rect 466 26901 522 26957
rect 590 26901 646 26957
rect 714 26901 770 26957
rect 838 26901 894 26957
rect 95 26440 151 26496
rect 219 26440 275 26496
rect 343 26440 399 26496
rect 467 26440 523 26496
rect 591 26440 647 26496
rect 715 26440 771 26496
rect 839 26440 895 26496
rect 95 26316 151 26372
rect 219 26316 275 26372
rect 343 26316 399 26372
rect 467 26316 523 26372
rect 591 26316 647 26372
rect 715 26316 771 26372
rect 839 26316 895 26372
rect 95 26192 151 26248
rect 219 26192 275 26248
rect 343 26192 399 26248
rect 467 26192 523 26248
rect 591 26192 647 26248
rect 715 26192 771 26248
rect 839 26192 895 26248
rect 95 26068 151 26124
rect 219 26068 275 26124
rect 343 26068 399 26124
rect 467 26068 523 26124
rect 591 26068 647 26124
rect 715 26068 771 26124
rect 839 26068 895 26124
rect 95 25944 151 26000
rect 219 25944 275 26000
rect 343 25944 399 26000
rect 467 25944 523 26000
rect 591 25944 647 26000
rect 715 25944 771 26000
rect 839 25944 895 26000
rect 95 25820 151 25876
rect 219 25820 275 25876
rect 343 25820 399 25876
rect 467 25820 523 25876
rect 591 25820 647 25876
rect 715 25820 771 25876
rect 839 25820 895 25876
rect 95 25696 151 25752
rect 219 25696 275 25752
rect 343 25696 399 25752
rect 467 25696 523 25752
rect 591 25696 647 25752
rect 715 25696 771 25752
rect 839 25696 895 25752
rect 95 25572 151 25628
rect 219 25572 275 25628
rect 343 25572 399 25628
rect 467 25572 523 25628
rect 591 25572 647 25628
rect 715 25572 771 25628
rect 839 25572 895 25628
rect 95 25448 151 25504
rect 219 25448 275 25504
rect 343 25448 399 25504
rect 467 25448 523 25504
rect 591 25448 647 25504
rect 715 25448 771 25504
rect 839 25448 895 25504
rect 95 25324 151 25380
rect 219 25324 275 25380
rect 343 25324 399 25380
rect 467 25324 523 25380
rect 591 25324 647 25380
rect 715 25324 771 25380
rect 839 25324 895 25380
rect 95 24828 151 24884
rect 219 24828 275 24884
rect 343 24828 399 24884
rect 467 24828 523 24884
rect 591 24828 647 24884
rect 715 24828 771 24884
rect 839 24828 895 24884
rect 95 24704 151 24760
rect 219 24704 275 24760
rect 343 24704 399 24760
rect 467 24704 523 24760
rect 591 24704 647 24760
rect 715 24704 771 24760
rect 839 24704 895 24760
rect 95 24580 151 24636
rect 219 24580 275 24636
rect 343 24580 399 24636
rect 467 24580 523 24636
rect 591 24580 647 24636
rect 715 24580 771 24636
rect 839 24580 895 24636
rect 95 24456 151 24512
rect 219 24456 275 24512
rect 343 24456 399 24512
rect 467 24456 523 24512
rect 591 24456 647 24512
rect 715 24456 771 24512
rect 839 24456 895 24512
rect 95 24332 151 24388
rect 219 24332 275 24388
rect 343 24332 399 24388
rect 467 24332 523 24388
rect 591 24332 647 24388
rect 715 24332 771 24388
rect 839 24332 895 24388
rect 95 24208 151 24264
rect 219 24208 275 24264
rect 343 24208 399 24264
rect 467 24208 523 24264
rect 591 24208 647 24264
rect 715 24208 771 24264
rect 839 24208 895 24264
rect 95 24084 151 24140
rect 219 24084 275 24140
rect 343 24084 399 24140
rect 467 24084 523 24140
rect 591 24084 647 24140
rect 715 24084 771 24140
rect 839 24084 895 24140
rect 95 23960 151 24016
rect 219 23960 275 24016
rect 343 23960 399 24016
rect 467 23960 523 24016
rect 591 23960 647 24016
rect 715 23960 771 24016
rect 839 23960 895 24016
rect 95 23836 151 23892
rect 219 23836 275 23892
rect 343 23836 399 23892
rect 467 23836 523 23892
rect 591 23836 647 23892
rect 715 23836 771 23892
rect 839 23836 895 23892
rect 95 23712 151 23768
rect 219 23712 275 23768
rect 343 23712 399 23768
rect 467 23712 523 23768
rect 591 23712 647 23768
rect 715 23712 771 23768
rect 839 23712 895 23768
rect 94 23241 150 23297
rect 218 23241 274 23297
rect 342 23241 398 23297
rect 466 23241 522 23297
rect 590 23241 646 23297
rect 714 23241 770 23297
rect 838 23241 894 23297
rect 94 23117 150 23173
rect 218 23117 274 23173
rect 342 23117 398 23173
rect 466 23117 522 23173
rect 590 23117 646 23173
rect 714 23117 770 23173
rect 838 23117 894 23173
rect 94 22993 150 23049
rect 218 22993 274 23049
rect 342 22993 398 23049
rect 466 22993 522 23049
rect 590 22993 646 23049
rect 714 22993 770 23049
rect 838 22993 894 23049
rect 94 22869 150 22925
rect 218 22869 274 22925
rect 342 22869 398 22925
rect 466 22869 522 22925
rect 590 22869 646 22925
rect 714 22869 770 22925
rect 838 22869 894 22925
rect 94 22745 150 22801
rect 218 22745 274 22801
rect 342 22745 398 22801
rect 466 22745 522 22801
rect 590 22745 646 22801
rect 714 22745 770 22801
rect 838 22745 894 22801
rect 94 22621 150 22677
rect 218 22621 274 22677
rect 342 22621 398 22677
rect 466 22621 522 22677
rect 590 22621 646 22677
rect 714 22621 770 22677
rect 838 22621 894 22677
rect 94 22497 150 22553
rect 218 22497 274 22553
rect 342 22497 398 22553
rect 466 22497 522 22553
rect 590 22497 646 22553
rect 714 22497 770 22553
rect 838 22497 894 22553
rect 94 22373 150 22429
rect 218 22373 274 22429
rect 342 22373 398 22429
rect 466 22373 522 22429
rect 590 22373 646 22429
rect 714 22373 770 22429
rect 838 22373 894 22429
rect 94 22249 150 22305
rect 218 22249 274 22305
rect 342 22249 398 22305
rect 466 22249 522 22305
rect 590 22249 646 22305
rect 714 22249 770 22305
rect 838 22249 894 22305
rect 94 22125 150 22181
rect 218 22125 274 22181
rect 342 22125 398 22181
rect 466 22125 522 22181
rect 590 22125 646 22181
rect 714 22125 770 22181
rect 838 22125 894 22181
rect 94 22001 150 22057
rect 218 22001 274 22057
rect 342 22001 398 22057
rect 466 22001 522 22057
rect 590 22001 646 22057
rect 714 22001 770 22057
rect 838 22001 894 22057
rect 94 21877 150 21933
rect 218 21877 274 21933
rect 342 21877 398 21933
rect 466 21877 522 21933
rect 590 21877 646 21933
rect 714 21877 770 21933
rect 838 21877 894 21933
rect 94 21753 150 21809
rect 218 21753 274 21809
rect 342 21753 398 21809
rect 466 21753 522 21809
rect 590 21753 646 21809
rect 714 21753 770 21809
rect 838 21753 894 21809
rect 94 21629 150 21685
rect 218 21629 274 21685
rect 342 21629 398 21685
rect 466 21629 522 21685
rect 590 21629 646 21685
rect 714 21629 770 21685
rect 838 21629 894 21685
rect 94 21505 150 21561
rect 218 21505 274 21561
rect 342 21505 398 21561
rect 466 21505 522 21561
rect 590 21505 646 21561
rect 714 21505 770 21561
rect 838 21505 894 21561
rect 94 21381 150 21437
rect 218 21381 274 21437
rect 342 21381 398 21437
rect 466 21381 522 21437
rect 590 21381 646 21437
rect 714 21381 770 21437
rect 838 21381 894 21437
rect 94 21257 150 21313
rect 218 21257 274 21313
rect 342 21257 398 21313
rect 466 21257 522 21313
rect 590 21257 646 21313
rect 714 21257 770 21313
rect 838 21257 894 21313
rect 94 21133 150 21189
rect 218 21133 274 21189
rect 342 21133 398 21189
rect 466 21133 522 21189
rect 590 21133 646 21189
rect 714 21133 770 21189
rect 838 21133 894 21189
rect 94 21009 150 21065
rect 218 21009 274 21065
rect 342 21009 398 21065
rect 466 21009 522 21065
rect 590 21009 646 21065
rect 714 21009 770 21065
rect 838 21009 894 21065
rect 94 20885 150 20941
rect 218 20885 274 20941
rect 342 20885 398 20941
rect 466 20885 522 20941
rect 590 20885 646 20941
rect 714 20885 770 20941
rect 838 20885 894 20941
rect 94 20761 150 20817
rect 218 20761 274 20817
rect 342 20761 398 20817
rect 466 20761 522 20817
rect 590 20761 646 20817
rect 714 20761 770 20817
rect 838 20761 894 20817
rect 94 20637 150 20693
rect 218 20637 274 20693
rect 342 20637 398 20693
rect 466 20637 522 20693
rect 590 20637 646 20693
rect 714 20637 770 20693
rect 838 20637 894 20693
rect 94 20513 150 20569
rect 218 20513 274 20569
rect 342 20513 398 20569
rect 466 20513 522 20569
rect 590 20513 646 20569
rect 714 20513 770 20569
rect 838 20513 894 20569
rect 94 20030 150 20086
rect 218 20030 274 20086
rect 342 20030 398 20086
rect 466 20030 522 20086
rect 590 20030 646 20086
rect 714 20030 770 20086
rect 838 20030 894 20086
rect 94 19906 150 19962
rect 218 19906 274 19962
rect 342 19906 398 19962
rect 466 19906 522 19962
rect 590 19906 646 19962
rect 714 19906 770 19962
rect 838 19906 894 19962
rect 94 19782 150 19838
rect 218 19782 274 19838
rect 342 19782 398 19838
rect 466 19782 522 19838
rect 590 19782 646 19838
rect 714 19782 770 19838
rect 838 19782 894 19838
rect 94 19658 150 19714
rect 218 19658 274 19714
rect 342 19658 398 19714
rect 466 19658 522 19714
rect 590 19658 646 19714
rect 714 19658 770 19714
rect 838 19658 894 19714
rect 94 19534 150 19590
rect 218 19534 274 19590
rect 342 19534 398 19590
rect 466 19534 522 19590
rect 590 19534 646 19590
rect 714 19534 770 19590
rect 838 19534 894 19590
rect 94 19410 150 19466
rect 218 19410 274 19466
rect 342 19410 398 19466
rect 466 19410 522 19466
rect 590 19410 646 19466
rect 714 19410 770 19466
rect 838 19410 894 19466
rect 94 19286 150 19342
rect 218 19286 274 19342
rect 342 19286 398 19342
rect 466 19286 522 19342
rect 590 19286 646 19342
rect 714 19286 770 19342
rect 838 19286 894 19342
rect 94 19162 150 19218
rect 218 19162 274 19218
rect 342 19162 398 19218
rect 466 19162 522 19218
rect 590 19162 646 19218
rect 714 19162 770 19218
rect 838 19162 894 19218
rect 94 19038 150 19094
rect 218 19038 274 19094
rect 342 19038 398 19094
rect 466 19038 522 19094
rect 590 19038 646 19094
rect 714 19038 770 19094
rect 838 19038 894 19094
rect 94 18914 150 18970
rect 218 18914 274 18970
rect 342 18914 398 18970
rect 466 18914 522 18970
rect 590 18914 646 18970
rect 714 18914 770 18970
rect 838 18914 894 18970
rect 94 18790 150 18846
rect 218 18790 274 18846
rect 342 18790 398 18846
rect 466 18790 522 18846
rect 590 18790 646 18846
rect 714 18790 770 18846
rect 838 18790 894 18846
rect 94 18666 150 18722
rect 218 18666 274 18722
rect 342 18666 398 18722
rect 466 18666 522 18722
rect 590 18666 646 18722
rect 714 18666 770 18722
rect 838 18666 894 18722
rect 94 18542 150 18598
rect 218 18542 274 18598
rect 342 18542 398 18598
rect 466 18542 522 18598
rect 590 18542 646 18598
rect 714 18542 770 18598
rect 838 18542 894 18598
rect 94 18418 150 18474
rect 218 18418 274 18474
rect 342 18418 398 18474
rect 466 18418 522 18474
rect 590 18418 646 18474
rect 714 18418 770 18474
rect 838 18418 894 18474
rect 94 18294 150 18350
rect 218 18294 274 18350
rect 342 18294 398 18350
rect 466 18294 522 18350
rect 590 18294 646 18350
rect 714 18294 770 18350
rect 838 18294 894 18350
rect 94 18170 150 18226
rect 218 18170 274 18226
rect 342 18170 398 18226
rect 466 18170 522 18226
rect 590 18170 646 18226
rect 714 18170 770 18226
rect 838 18170 894 18226
rect 94 18046 150 18102
rect 218 18046 274 18102
rect 342 18046 398 18102
rect 466 18046 522 18102
rect 590 18046 646 18102
rect 714 18046 770 18102
rect 838 18046 894 18102
rect 94 17922 150 17978
rect 218 17922 274 17978
rect 342 17922 398 17978
rect 466 17922 522 17978
rect 590 17922 646 17978
rect 714 17922 770 17978
rect 838 17922 894 17978
rect 94 17798 150 17854
rect 218 17798 274 17854
rect 342 17798 398 17854
rect 466 17798 522 17854
rect 590 17798 646 17854
rect 714 17798 770 17854
rect 838 17798 894 17854
rect 94 17674 150 17730
rect 218 17674 274 17730
rect 342 17674 398 17730
rect 466 17674 522 17730
rect 590 17674 646 17730
rect 714 17674 770 17730
rect 838 17674 894 17730
rect 94 17550 150 17606
rect 218 17550 274 17606
rect 342 17550 398 17606
rect 466 17550 522 17606
rect 590 17550 646 17606
rect 714 17550 770 17606
rect 838 17550 894 17606
rect 94 17426 150 17482
rect 218 17426 274 17482
rect 342 17426 398 17482
rect 466 17426 522 17482
rect 590 17426 646 17482
rect 714 17426 770 17482
rect 838 17426 894 17482
rect 94 17302 150 17358
rect 218 17302 274 17358
rect 342 17302 398 17358
rect 466 17302 522 17358
rect 590 17302 646 17358
rect 714 17302 770 17358
rect 838 17302 894 17358
rect 94 16857 150 16913
rect 218 16857 274 16913
rect 342 16857 398 16913
rect 466 16857 522 16913
rect 590 16857 646 16913
rect 714 16857 770 16913
rect 838 16857 894 16913
rect 94 16733 150 16789
rect 218 16733 274 16789
rect 342 16733 398 16789
rect 466 16733 522 16789
rect 590 16733 646 16789
rect 714 16733 770 16789
rect 838 16733 894 16789
rect 94 16609 150 16665
rect 218 16609 274 16665
rect 342 16609 398 16665
rect 466 16609 522 16665
rect 590 16609 646 16665
rect 714 16609 770 16665
rect 838 16609 894 16665
rect 94 16485 150 16541
rect 218 16485 274 16541
rect 342 16485 398 16541
rect 466 16485 522 16541
rect 590 16485 646 16541
rect 714 16485 770 16541
rect 838 16485 894 16541
rect 94 16361 150 16417
rect 218 16361 274 16417
rect 342 16361 398 16417
rect 466 16361 522 16417
rect 590 16361 646 16417
rect 714 16361 770 16417
rect 838 16361 894 16417
rect 94 16237 150 16293
rect 218 16237 274 16293
rect 342 16237 398 16293
rect 466 16237 522 16293
rect 590 16237 646 16293
rect 714 16237 770 16293
rect 838 16237 894 16293
rect 94 16113 150 16169
rect 218 16113 274 16169
rect 342 16113 398 16169
rect 466 16113 522 16169
rect 590 16113 646 16169
rect 714 16113 770 16169
rect 838 16113 894 16169
rect 94 15989 150 16045
rect 218 15989 274 16045
rect 342 15989 398 16045
rect 466 15989 522 16045
rect 590 15989 646 16045
rect 714 15989 770 16045
rect 838 15989 894 16045
rect 94 15865 150 15921
rect 218 15865 274 15921
rect 342 15865 398 15921
rect 466 15865 522 15921
rect 590 15865 646 15921
rect 714 15865 770 15921
rect 838 15865 894 15921
rect 94 15741 150 15797
rect 218 15741 274 15797
rect 342 15741 398 15797
rect 466 15741 522 15797
rect 590 15741 646 15797
rect 714 15741 770 15797
rect 838 15741 894 15797
rect 94 15617 150 15673
rect 218 15617 274 15673
rect 342 15617 398 15673
rect 466 15617 522 15673
rect 590 15617 646 15673
rect 714 15617 770 15673
rect 838 15617 894 15673
rect 94 15493 150 15549
rect 218 15493 274 15549
rect 342 15493 398 15549
rect 466 15493 522 15549
rect 590 15493 646 15549
rect 714 15493 770 15549
rect 838 15493 894 15549
rect 94 15369 150 15425
rect 218 15369 274 15425
rect 342 15369 398 15425
rect 466 15369 522 15425
rect 590 15369 646 15425
rect 714 15369 770 15425
rect 838 15369 894 15425
rect 94 15245 150 15301
rect 218 15245 274 15301
rect 342 15245 398 15301
rect 466 15245 522 15301
rect 590 15245 646 15301
rect 714 15245 770 15301
rect 838 15245 894 15301
rect 94 15121 150 15177
rect 218 15121 274 15177
rect 342 15121 398 15177
rect 466 15121 522 15177
rect 590 15121 646 15177
rect 714 15121 770 15177
rect 838 15121 894 15177
rect 94 14997 150 15053
rect 218 14997 274 15053
rect 342 14997 398 15053
rect 466 14997 522 15053
rect 590 14997 646 15053
rect 714 14997 770 15053
rect 838 14997 894 15053
rect 94 14873 150 14929
rect 218 14873 274 14929
rect 342 14873 398 14929
rect 466 14873 522 14929
rect 590 14873 646 14929
rect 714 14873 770 14929
rect 838 14873 894 14929
rect 94 14749 150 14805
rect 218 14749 274 14805
rect 342 14749 398 14805
rect 466 14749 522 14805
rect 590 14749 646 14805
rect 714 14749 770 14805
rect 838 14749 894 14805
rect 94 14625 150 14681
rect 218 14625 274 14681
rect 342 14625 398 14681
rect 466 14625 522 14681
rect 590 14625 646 14681
rect 714 14625 770 14681
rect 838 14625 894 14681
rect 94 14501 150 14557
rect 218 14501 274 14557
rect 342 14501 398 14557
rect 466 14501 522 14557
rect 590 14501 646 14557
rect 714 14501 770 14557
rect 838 14501 894 14557
rect 94 14377 150 14433
rect 218 14377 274 14433
rect 342 14377 398 14433
rect 466 14377 522 14433
rect 590 14377 646 14433
rect 714 14377 770 14433
rect 838 14377 894 14433
rect 94 14253 150 14309
rect 218 14253 274 14309
rect 342 14253 398 14309
rect 466 14253 522 14309
rect 590 14253 646 14309
rect 714 14253 770 14309
rect 838 14253 894 14309
rect 94 14129 150 14185
rect 218 14129 274 14185
rect 342 14129 398 14185
rect 466 14129 522 14185
rect 590 14129 646 14185
rect 714 14129 770 14185
rect 838 14129 894 14185
<< metal4 >>
rect 0 69629 1000 69678
rect 0 69573 94 69629
rect 150 69573 218 69629
rect 274 69573 342 69629
rect 398 69573 466 69629
rect 522 69573 590 69629
rect 646 69573 714 69629
rect 770 69573 838 69629
rect 894 69573 1000 69629
rect 0 69505 1000 69573
rect 0 69449 94 69505
rect 150 69449 218 69505
rect 274 69449 342 69505
rect 398 69449 466 69505
rect 522 69449 590 69505
rect 646 69449 714 69505
rect 770 69449 838 69505
rect 894 69449 1000 69505
rect 0 69381 1000 69449
rect 0 69325 94 69381
rect 150 69325 218 69381
rect 274 69325 342 69381
rect 398 69325 466 69381
rect 522 69325 590 69381
rect 646 69325 714 69381
rect 770 69325 838 69381
rect 894 69325 1000 69381
rect 0 69257 1000 69325
rect 0 69201 94 69257
rect 150 69201 218 69257
rect 274 69201 342 69257
rect 398 69201 466 69257
rect 522 69201 590 69257
rect 646 69201 714 69257
rect 770 69201 838 69257
rect 894 69201 1000 69257
rect 0 69133 1000 69201
rect 0 69077 94 69133
rect 150 69077 218 69133
rect 274 69077 342 69133
rect 398 69077 466 69133
rect 522 69077 590 69133
rect 646 69077 714 69133
rect 770 69077 838 69133
rect 894 69077 1000 69133
rect 0 69009 1000 69077
rect 0 68953 94 69009
rect 150 68953 218 69009
rect 274 68953 342 69009
rect 398 68953 466 69009
rect 522 68953 590 69009
rect 646 68953 714 69009
rect 770 68953 838 69009
rect 894 68953 1000 69009
rect 0 68885 1000 68953
rect 0 68829 94 68885
rect 150 68829 218 68885
rect 274 68829 342 68885
rect 398 68829 466 68885
rect 522 68829 590 68885
rect 646 68829 714 68885
rect 770 68829 838 68885
rect 894 68829 1000 68885
rect 0 68761 1000 68829
rect 0 68705 94 68761
rect 150 68705 218 68761
rect 274 68705 342 68761
rect 398 68705 466 68761
rect 522 68705 590 68761
rect 646 68705 714 68761
rect 770 68705 838 68761
rect 894 68705 1000 68761
rect 0 68637 1000 68705
rect 0 68581 94 68637
rect 150 68581 218 68637
rect 274 68581 342 68637
rect 398 68581 466 68637
rect 522 68581 590 68637
rect 646 68581 714 68637
rect 770 68581 838 68637
rect 894 68581 1000 68637
rect 0 68513 1000 68581
rect 0 68457 94 68513
rect 150 68457 218 68513
rect 274 68457 342 68513
rect 398 68457 466 68513
rect 522 68457 590 68513
rect 646 68457 714 68513
rect 770 68457 838 68513
rect 894 68457 1000 68513
rect 0 68400 1000 68457
rect 0 68084 1000 68200
rect 0 68028 94 68084
rect 150 68028 218 68084
rect 274 68028 342 68084
rect 398 68028 466 68084
rect 522 68028 590 68084
rect 646 68028 714 68084
rect 770 68028 838 68084
rect 894 68028 1000 68084
rect 0 67960 1000 68028
rect 0 67904 94 67960
rect 150 67904 218 67960
rect 274 67904 342 67960
rect 398 67904 466 67960
rect 522 67904 590 67960
rect 646 67904 714 67960
rect 770 67904 838 67960
rect 894 67904 1000 67960
rect 0 67836 1000 67904
rect 0 67780 94 67836
rect 150 67780 218 67836
rect 274 67780 342 67836
rect 398 67780 466 67836
rect 522 67780 590 67836
rect 646 67780 714 67836
rect 770 67780 838 67836
rect 894 67780 1000 67836
rect 0 67712 1000 67780
rect 0 67656 94 67712
rect 150 67656 218 67712
rect 274 67656 342 67712
rect 398 67656 466 67712
rect 522 67656 590 67712
rect 646 67656 714 67712
rect 770 67656 838 67712
rect 894 67656 1000 67712
rect 0 67588 1000 67656
rect 0 67532 94 67588
rect 150 67532 218 67588
rect 274 67532 342 67588
rect 398 67532 466 67588
rect 522 67532 590 67588
rect 646 67532 714 67588
rect 770 67532 838 67588
rect 894 67532 1000 67588
rect 0 67464 1000 67532
rect 0 67408 94 67464
rect 150 67408 218 67464
rect 274 67408 342 67464
rect 398 67408 466 67464
rect 522 67408 590 67464
rect 646 67408 714 67464
rect 770 67408 838 67464
rect 894 67408 1000 67464
rect 0 67340 1000 67408
rect 0 67284 94 67340
rect 150 67284 218 67340
rect 274 67284 342 67340
rect 398 67284 466 67340
rect 522 67284 590 67340
rect 646 67284 714 67340
rect 770 67284 838 67340
rect 894 67284 1000 67340
rect 0 67216 1000 67284
rect 0 67160 94 67216
rect 150 67160 218 67216
rect 274 67160 342 67216
rect 398 67160 466 67216
rect 522 67160 590 67216
rect 646 67160 714 67216
rect 770 67160 838 67216
rect 894 67160 1000 67216
rect 0 67092 1000 67160
rect 0 67036 94 67092
rect 150 67036 218 67092
rect 274 67036 342 67092
rect 398 67036 466 67092
rect 522 67036 590 67092
rect 646 67036 714 67092
rect 770 67036 838 67092
rect 894 67036 1000 67092
rect 0 66968 1000 67036
rect 0 66912 94 66968
rect 150 66912 218 66968
rect 274 66912 342 66968
rect 398 66912 466 66968
rect 522 66912 590 66968
rect 646 66912 714 66968
rect 770 66912 838 66968
rect 894 66912 1000 66968
rect 0 66800 1000 66912
rect 0 66477 1000 66600
rect 0 66421 94 66477
rect 150 66421 218 66477
rect 274 66421 342 66477
rect 398 66421 466 66477
rect 522 66421 590 66477
rect 646 66421 714 66477
rect 770 66421 838 66477
rect 894 66421 1000 66477
rect 0 66353 1000 66421
rect 0 66297 94 66353
rect 150 66297 218 66353
rect 274 66297 342 66353
rect 398 66297 466 66353
rect 522 66297 590 66353
rect 646 66297 714 66353
rect 770 66297 838 66353
rect 894 66297 1000 66353
rect 0 66229 1000 66297
rect 0 66173 94 66229
rect 150 66173 218 66229
rect 274 66173 342 66229
rect 398 66173 466 66229
rect 522 66173 590 66229
rect 646 66173 714 66229
rect 770 66173 838 66229
rect 894 66173 1000 66229
rect 0 66105 1000 66173
rect 0 66049 94 66105
rect 150 66049 218 66105
rect 274 66049 342 66105
rect 398 66049 466 66105
rect 522 66049 590 66105
rect 646 66049 714 66105
rect 770 66049 838 66105
rect 894 66049 1000 66105
rect 0 65981 1000 66049
rect 0 65925 94 65981
rect 150 65925 218 65981
rect 274 65925 342 65981
rect 398 65925 466 65981
rect 522 65925 590 65981
rect 646 65925 714 65981
rect 770 65925 838 65981
rect 894 65925 1000 65981
rect 0 65857 1000 65925
rect 0 65801 94 65857
rect 150 65801 218 65857
rect 274 65801 342 65857
rect 398 65801 466 65857
rect 522 65801 590 65857
rect 646 65801 714 65857
rect 770 65801 838 65857
rect 894 65801 1000 65857
rect 0 65733 1000 65801
rect 0 65677 94 65733
rect 150 65677 218 65733
rect 274 65677 342 65733
rect 398 65677 466 65733
rect 522 65677 590 65733
rect 646 65677 714 65733
rect 770 65677 838 65733
rect 894 65677 1000 65733
rect 0 65609 1000 65677
rect 0 65553 94 65609
rect 150 65553 218 65609
rect 274 65553 342 65609
rect 398 65553 466 65609
rect 522 65553 590 65609
rect 646 65553 714 65609
rect 770 65553 838 65609
rect 894 65553 1000 65609
rect 0 65485 1000 65553
rect 0 65429 94 65485
rect 150 65429 218 65485
rect 274 65429 342 65485
rect 398 65429 466 65485
rect 522 65429 590 65485
rect 646 65429 714 65485
rect 770 65429 838 65485
rect 894 65429 1000 65485
rect 0 65361 1000 65429
rect 0 65305 94 65361
rect 150 65305 218 65361
rect 274 65305 342 65361
rect 398 65305 466 65361
rect 522 65305 590 65361
rect 646 65305 714 65361
rect 770 65305 838 65361
rect 894 65305 1000 65361
rect 0 65200 1000 65305
rect 0 64886 1000 65000
rect 0 64830 94 64886
rect 150 64830 218 64886
rect 274 64830 342 64886
rect 398 64830 466 64886
rect 522 64830 590 64886
rect 646 64830 714 64886
rect 770 64830 838 64886
rect 894 64830 1000 64886
rect 0 64762 1000 64830
rect 0 64706 94 64762
rect 150 64706 218 64762
rect 274 64706 342 64762
rect 398 64706 466 64762
rect 522 64706 590 64762
rect 646 64706 714 64762
rect 770 64706 838 64762
rect 894 64706 1000 64762
rect 0 64638 1000 64706
rect 0 64582 94 64638
rect 150 64582 218 64638
rect 274 64582 342 64638
rect 398 64582 466 64638
rect 522 64582 590 64638
rect 646 64582 714 64638
rect 770 64582 838 64638
rect 894 64582 1000 64638
rect 0 64514 1000 64582
rect 0 64458 94 64514
rect 150 64458 218 64514
rect 274 64458 342 64514
rect 398 64458 466 64514
rect 522 64458 590 64514
rect 646 64458 714 64514
rect 770 64458 838 64514
rect 894 64458 1000 64514
rect 0 64390 1000 64458
rect 0 64334 94 64390
rect 150 64334 218 64390
rect 274 64334 342 64390
rect 398 64334 466 64390
rect 522 64334 590 64390
rect 646 64334 714 64390
rect 770 64334 838 64390
rect 894 64334 1000 64390
rect 0 64266 1000 64334
rect 0 64210 94 64266
rect 150 64210 218 64266
rect 274 64210 342 64266
rect 398 64210 466 64266
rect 522 64210 590 64266
rect 646 64210 714 64266
rect 770 64210 838 64266
rect 894 64210 1000 64266
rect 0 64142 1000 64210
rect 0 64086 94 64142
rect 150 64086 218 64142
rect 274 64086 342 64142
rect 398 64086 466 64142
rect 522 64086 590 64142
rect 646 64086 714 64142
rect 770 64086 838 64142
rect 894 64086 1000 64142
rect 0 64018 1000 64086
rect 0 63962 94 64018
rect 150 63962 218 64018
rect 274 63962 342 64018
rect 398 63962 466 64018
rect 522 63962 590 64018
rect 646 63962 714 64018
rect 770 63962 838 64018
rect 894 63962 1000 64018
rect 0 63894 1000 63962
rect 0 63838 94 63894
rect 150 63838 218 63894
rect 274 63838 342 63894
rect 398 63838 466 63894
rect 522 63838 590 63894
rect 646 63838 714 63894
rect 770 63838 838 63894
rect 894 63838 1000 63894
rect 0 63770 1000 63838
rect 0 63714 94 63770
rect 150 63714 218 63770
rect 274 63714 342 63770
rect 398 63714 466 63770
rect 522 63714 590 63770
rect 646 63714 714 63770
rect 770 63714 838 63770
rect 894 63714 1000 63770
rect 0 63600 1000 63714
rect 0 63280 1000 63400
rect 0 63224 94 63280
rect 150 63224 218 63280
rect 274 63224 342 63280
rect 398 63224 466 63280
rect 522 63224 590 63280
rect 646 63224 714 63280
rect 770 63224 838 63280
rect 894 63224 1000 63280
rect 0 63156 1000 63224
rect 0 63100 94 63156
rect 150 63100 218 63156
rect 274 63100 342 63156
rect 398 63100 466 63156
rect 522 63100 590 63156
rect 646 63100 714 63156
rect 770 63100 838 63156
rect 894 63100 1000 63156
rect 0 63032 1000 63100
rect 0 62976 94 63032
rect 150 62976 218 63032
rect 274 62976 342 63032
rect 398 62976 466 63032
rect 522 62976 590 63032
rect 646 62976 714 63032
rect 770 62976 838 63032
rect 894 62976 1000 63032
rect 0 62908 1000 62976
rect 0 62852 94 62908
rect 150 62852 218 62908
rect 274 62852 342 62908
rect 398 62852 466 62908
rect 522 62852 590 62908
rect 646 62852 714 62908
rect 770 62852 838 62908
rect 894 62852 1000 62908
rect 0 62784 1000 62852
rect 0 62728 94 62784
rect 150 62728 218 62784
rect 274 62728 342 62784
rect 398 62728 466 62784
rect 522 62728 590 62784
rect 646 62728 714 62784
rect 770 62728 838 62784
rect 894 62728 1000 62784
rect 0 62660 1000 62728
rect 0 62604 94 62660
rect 150 62604 218 62660
rect 274 62604 342 62660
rect 398 62604 466 62660
rect 522 62604 590 62660
rect 646 62604 714 62660
rect 770 62604 838 62660
rect 894 62604 1000 62660
rect 0 62536 1000 62604
rect 0 62480 94 62536
rect 150 62480 218 62536
rect 274 62480 342 62536
rect 398 62480 466 62536
rect 522 62480 590 62536
rect 646 62480 714 62536
rect 770 62480 838 62536
rect 894 62480 1000 62536
rect 0 62412 1000 62480
rect 0 62356 94 62412
rect 150 62356 218 62412
rect 274 62356 342 62412
rect 398 62356 466 62412
rect 522 62356 590 62412
rect 646 62356 714 62412
rect 770 62356 838 62412
rect 894 62356 1000 62412
rect 0 62288 1000 62356
rect 0 62232 94 62288
rect 150 62232 218 62288
rect 274 62232 342 62288
rect 398 62232 466 62288
rect 522 62232 590 62288
rect 646 62232 714 62288
rect 770 62232 838 62288
rect 894 62232 1000 62288
rect 0 62164 1000 62232
rect 0 62108 94 62164
rect 150 62108 218 62164
rect 274 62108 342 62164
rect 398 62108 466 62164
rect 522 62108 590 62164
rect 646 62108 714 62164
rect 770 62108 838 62164
rect 894 62108 1000 62164
rect 0 62000 1000 62108
rect 0 61694 1000 61800
rect 0 61638 94 61694
rect 150 61638 218 61694
rect 274 61638 342 61694
rect 398 61638 466 61694
rect 522 61638 590 61694
rect 646 61638 714 61694
rect 770 61638 838 61694
rect 894 61638 1000 61694
rect 0 61570 1000 61638
rect 0 61514 94 61570
rect 150 61514 218 61570
rect 274 61514 342 61570
rect 398 61514 466 61570
rect 522 61514 590 61570
rect 646 61514 714 61570
rect 770 61514 838 61570
rect 894 61514 1000 61570
rect 0 61446 1000 61514
rect 0 61390 94 61446
rect 150 61390 218 61446
rect 274 61390 342 61446
rect 398 61390 466 61446
rect 522 61390 590 61446
rect 646 61390 714 61446
rect 770 61390 838 61446
rect 894 61390 1000 61446
rect 0 61322 1000 61390
rect 0 61266 94 61322
rect 150 61266 218 61322
rect 274 61266 342 61322
rect 398 61266 466 61322
rect 522 61266 590 61322
rect 646 61266 714 61322
rect 770 61266 838 61322
rect 894 61266 1000 61322
rect 0 61198 1000 61266
rect 0 61142 94 61198
rect 150 61142 218 61198
rect 274 61142 342 61198
rect 398 61142 466 61198
rect 522 61142 590 61198
rect 646 61142 714 61198
rect 770 61142 838 61198
rect 894 61142 1000 61198
rect 0 61074 1000 61142
rect 0 61018 94 61074
rect 150 61018 218 61074
rect 274 61018 342 61074
rect 398 61018 466 61074
rect 522 61018 590 61074
rect 646 61018 714 61074
rect 770 61018 838 61074
rect 894 61018 1000 61074
rect 0 60950 1000 61018
rect 0 60894 94 60950
rect 150 60894 218 60950
rect 274 60894 342 60950
rect 398 60894 466 60950
rect 522 60894 590 60950
rect 646 60894 714 60950
rect 770 60894 838 60950
rect 894 60894 1000 60950
rect 0 60826 1000 60894
rect 0 60770 94 60826
rect 150 60770 218 60826
rect 274 60770 342 60826
rect 398 60770 466 60826
rect 522 60770 590 60826
rect 646 60770 714 60826
rect 770 60770 838 60826
rect 894 60770 1000 60826
rect 0 60702 1000 60770
rect 0 60646 94 60702
rect 150 60646 218 60702
rect 274 60646 342 60702
rect 398 60646 466 60702
rect 522 60646 590 60702
rect 646 60646 714 60702
rect 770 60646 838 60702
rect 894 60646 1000 60702
rect 0 60578 1000 60646
rect 0 60522 94 60578
rect 150 60522 218 60578
rect 274 60522 342 60578
rect 398 60522 466 60578
rect 522 60522 590 60578
rect 646 60522 714 60578
rect 770 60522 838 60578
rect 894 60522 1000 60578
rect 0 60400 1000 60522
rect 0 60102 1000 60200
rect 0 60046 94 60102
rect 150 60046 218 60102
rect 274 60046 342 60102
rect 398 60046 466 60102
rect 522 60046 590 60102
rect 646 60046 714 60102
rect 770 60046 838 60102
rect 894 60046 1000 60102
rect 0 59978 1000 60046
rect 0 59922 94 59978
rect 150 59922 218 59978
rect 274 59922 342 59978
rect 398 59922 466 59978
rect 522 59922 590 59978
rect 646 59922 714 59978
rect 770 59922 838 59978
rect 894 59922 1000 59978
rect 0 59854 1000 59922
rect 0 59798 94 59854
rect 150 59798 218 59854
rect 274 59798 342 59854
rect 398 59798 466 59854
rect 522 59798 590 59854
rect 646 59798 714 59854
rect 770 59798 838 59854
rect 894 59798 1000 59854
rect 0 59730 1000 59798
rect 0 59674 94 59730
rect 150 59674 218 59730
rect 274 59674 342 59730
rect 398 59674 466 59730
rect 522 59674 590 59730
rect 646 59674 714 59730
rect 770 59674 838 59730
rect 894 59674 1000 59730
rect 0 59606 1000 59674
rect 0 59550 94 59606
rect 150 59550 218 59606
rect 274 59550 342 59606
rect 398 59550 466 59606
rect 522 59550 590 59606
rect 646 59550 714 59606
rect 770 59550 838 59606
rect 894 59550 1000 59606
rect 0 59482 1000 59550
rect 0 59426 94 59482
rect 150 59426 218 59482
rect 274 59426 342 59482
rect 398 59426 466 59482
rect 522 59426 590 59482
rect 646 59426 714 59482
rect 770 59426 838 59482
rect 894 59426 1000 59482
rect 0 59358 1000 59426
rect 0 59302 94 59358
rect 150 59302 218 59358
rect 274 59302 342 59358
rect 398 59302 466 59358
rect 522 59302 590 59358
rect 646 59302 714 59358
rect 770 59302 838 59358
rect 894 59302 1000 59358
rect 0 59234 1000 59302
rect 0 59178 94 59234
rect 150 59178 218 59234
rect 274 59178 342 59234
rect 398 59178 466 59234
rect 522 59178 590 59234
rect 646 59178 714 59234
rect 770 59178 838 59234
rect 894 59178 1000 59234
rect 0 59110 1000 59178
rect 0 59054 94 59110
rect 150 59054 218 59110
rect 274 59054 342 59110
rect 398 59054 466 59110
rect 522 59054 590 59110
rect 646 59054 714 59110
rect 770 59054 838 59110
rect 894 59054 1000 59110
rect 0 58986 1000 59054
rect 0 58930 94 58986
rect 150 58930 218 58986
rect 274 58930 342 58986
rect 398 58930 466 58986
rect 522 58930 590 58986
rect 646 58930 714 58986
rect 770 58930 838 58986
rect 894 58930 1000 58986
rect 0 58800 1000 58930
rect 0 58485 1000 58600
rect 0 58429 94 58485
rect 150 58429 218 58485
rect 274 58429 342 58485
rect 398 58429 466 58485
rect 522 58429 590 58485
rect 646 58429 714 58485
rect 770 58429 838 58485
rect 894 58429 1000 58485
rect 0 58361 1000 58429
rect 0 58305 94 58361
rect 150 58305 218 58361
rect 274 58305 342 58361
rect 398 58305 466 58361
rect 522 58305 590 58361
rect 646 58305 714 58361
rect 770 58305 838 58361
rect 894 58305 1000 58361
rect 0 58237 1000 58305
rect 0 58181 94 58237
rect 150 58181 218 58237
rect 274 58181 342 58237
rect 398 58181 466 58237
rect 522 58181 590 58237
rect 646 58181 714 58237
rect 770 58181 838 58237
rect 894 58181 1000 58237
rect 0 58113 1000 58181
rect 0 58057 94 58113
rect 150 58057 218 58113
rect 274 58057 342 58113
rect 398 58057 466 58113
rect 522 58057 590 58113
rect 646 58057 714 58113
rect 770 58057 838 58113
rect 894 58057 1000 58113
rect 0 57989 1000 58057
rect 0 57933 94 57989
rect 150 57933 218 57989
rect 274 57933 342 57989
rect 398 57933 466 57989
rect 522 57933 590 57989
rect 646 57933 714 57989
rect 770 57933 838 57989
rect 894 57933 1000 57989
rect 0 57865 1000 57933
rect 0 57809 94 57865
rect 150 57809 218 57865
rect 274 57809 342 57865
rect 398 57809 466 57865
rect 522 57809 590 57865
rect 646 57809 714 57865
rect 770 57809 838 57865
rect 894 57809 1000 57865
rect 0 57741 1000 57809
rect 0 57685 94 57741
rect 150 57685 218 57741
rect 274 57685 342 57741
rect 398 57685 466 57741
rect 522 57685 590 57741
rect 646 57685 714 57741
rect 770 57685 838 57741
rect 894 57685 1000 57741
rect 0 57617 1000 57685
rect 0 57561 94 57617
rect 150 57561 218 57617
rect 274 57561 342 57617
rect 398 57561 466 57617
rect 522 57561 590 57617
rect 646 57561 714 57617
rect 770 57561 838 57617
rect 894 57561 1000 57617
rect 0 57493 1000 57561
rect 0 57437 94 57493
rect 150 57437 218 57493
rect 274 57437 342 57493
rect 398 57437 466 57493
rect 522 57437 590 57493
rect 646 57437 714 57493
rect 770 57437 838 57493
rect 894 57437 1000 57493
rect 0 57369 1000 57437
rect 0 57313 94 57369
rect 150 57313 218 57369
rect 274 57313 342 57369
rect 398 57313 466 57369
rect 522 57313 590 57369
rect 646 57313 714 57369
rect 770 57313 838 57369
rect 894 57313 1000 57369
rect 0 57200 1000 57313
rect 0 56892 1000 57000
rect 0 56836 94 56892
rect 150 56836 218 56892
rect 274 56836 342 56892
rect 398 56836 466 56892
rect 522 56836 590 56892
rect 646 56836 714 56892
rect 770 56836 838 56892
rect 894 56836 1000 56892
rect 0 56768 1000 56836
rect 0 56712 94 56768
rect 150 56712 218 56768
rect 274 56712 342 56768
rect 398 56712 466 56768
rect 522 56712 590 56768
rect 646 56712 714 56768
rect 770 56712 838 56768
rect 894 56712 1000 56768
rect 0 56644 1000 56712
rect 0 56588 94 56644
rect 150 56588 218 56644
rect 274 56588 342 56644
rect 398 56588 466 56644
rect 522 56588 590 56644
rect 646 56588 714 56644
rect 770 56588 838 56644
rect 894 56588 1000 56644
rect 0 56520 1000 56588
rect 0 56464 94 56520
rect 150 56464 218 56520
rect 274 56464 342 56520
rect 398 56464 466 56520
rect 522 56464 590 56520
rect 646 56464 714 56520
rect 770 56464 838 56520
rect 894 56464 1000 56520
rect 0 56396 1000 56464
rect 0 56340 94 56396
rect 150 56340 218 56396
rect 274 56340 342 56396
rect 398 56340 466 56396
rect 522 56340 590 56396
rect 646 56340 714 56396
rect 770 56340 838 56396
rect 894 56340 1000 56396
rect 0 56272 1000 56340
rect 0 56216 94 56272
rect 150 56216 218 56272
rect 274 56216 342 56272
rect 398 56216 466 56272
rect 522 56216 590 56272
rect 646 56216 714 56272
rect 770 56216 838 56272
rect 894 56216 1000 56272
rect 0 56148 1000 56216
rect 0 56092 94 56148
rect 150 56092 218 56148
rect 274 56092 342 56148
rect 398 56092 466 56148
rect 522 56092 590 56148
rect 646 56092 714 56148
rect 770 56092 838 56148
rect 894 56092 1000 56148
rect 0 56024 1000 56092
rect 0 55968 94 56024
rect 150 55968 218 56024
rect 274 55968 342 56024
rect 398 55968 466 56024
rect 522 55968 590 56024
rect 646 55968 714 56024
rect 770 55968 838 56024
rect 894 55968 1000 56024
rect 0 55900 1000 55968
rect 0 55844 94 55900
rect 150 55844 218 55900
rect 274 55844 342 55900
rect 398 55844 466 55900
rect 522 55844 590 55900
rect 646 55844 714 55900
rect 770 55844 838 55900
rect 894 55844 1000 55900
rect 0 55776 1000 55844
rect 0 55720 94 55776
rect 150 55720 218 55776
rect 274 55720 342 55776
rect 398 55720 466 55776
rect 522 55720 590 55776
rect 646 55720 714 55776
rect 770 55720 838 55776
rect 894 55720 1000 55776
rect 0 55600 1000 55720
rect 0 55288 1000 55400
rect 0 55232 94 55288
rect 150 55232 218 55288
rect 274 55232 342 55288
rect 398 55232 466 55288
rect 522 55232 590 55288
rect 646 55232 714 55288
rect 770 55232 838 55288
rect 894 55232 1000 55288
rect 0 55164 1000 55232
rect 0 55108 94 55164
rect 150 55108 218 55164
rect 274 55108 342 55164
rect 398 55108 466 55164
rect 522 55108 590 55164
rect 646 55108 714 55164
rect 770 55108 838 55164
rect 894 55108 1000 55164
rect 0 55040 1000 55108
rect 0 54984 94 55040
rect 150 54984 218 55040
rect 274 54984 342 55040
rect 398 54984 466 55040
rect 522 54984 590 55040
rect 646 54984 714 55040
rect 770 54984 838 55040
rect 894 54984 1000 55040
rect 0 54916 1000 54984
rect 0 54860 94 54916
rect 150 54860 218 54916
rect 274 54860 342 54916
rect 398 54860 466 54916
rect 522 54860 590 54916
rect 646 54860 714 54916
rect 770 54860 838 54916
rect 894 54860 1000 54916
rect 0 54792 1000 54860
rect 0 54736 94 54792
rect 150 54736 218 54792
rect 274 54736 342 54792
rect 398 54736 466 54792
rect 522 54736 590 54792
rect 646 54736 714 54792
rect 770 54736 838 54792
rect 894 54736 1000 54792
rect 0 54668 1000 54736
rect 0 54612 94 54668
rect 150 54612 218 54668
rect 274 54612 342 54668
rect 398 54612 466 54668
rect 522 54612 590 54668
rect 646 54612 714 54668
rect 770 54612 838 54668
rect 894 54612 1000 54668
rect 0 54544 1000 54612
rect 0 54488 94 54544
rect 150 54488 218 54544
rect 274 54488 342 54544
rect 398 54488 466 54544
rect 522 54488 590 54544
rect 646 54488 714 54544
rect 770 54488 838 54544
rect 894 54488 1000 54544
rect 0 54420 1000 54488
rect 0 54364 94 54420
rect 150 54364 218 54420
rect 274 54364 342 54420
rect 398 54364 466 54420
rect 522 54364 590 54420
rect 646 54364 714 54420
rect 770 54364 838 54420
rect 894 54364 1000 54420
rect 0 54296 1000 54364
rect 0 54240 94 54296
rect 150 54240 218 54296
rect 274 54240 342 54296
rect 398 54240 466 54296
rect 522 54240 590 54296
rect 646 54240 714 54296
rect 770 54240 838 54296
rect 894 54240 1000 54296
rect 0 54172 1000 54240
rect 0 54116 94 54172
rect 150 54116 218 54172
rect 274 54116 342 54172
rect 398 54116 466 54172
rect 522 54116 590 54172
rect 646 54116 714 54172
rect 770 54116 838 54172
rect 894 54116 1000 54172
rect 0 54000 1000 54116
rect 0 53682 1000 53800
rect 0 53626 94 53682
rect 150 53626 218 53682
rect 274 53626 342 53682
rect 398 53626 466 53682
rect 522 53626 590 53682
rect 646 53626 714 53682
rect 770 53626 838 53682
rect 894 53626 1000 53682
rect 0 53558 1000 53626
rect 0 53502 94 53558
rect 150 53502 218 53558
rect 274 53502 342 53558
rect 398 53502 466 53558
rect 522 53502 590 53558
rect 646 53502 714 53558
rect 770 53502 838 53558
rect 894 53502 1000 53558
rect 0 53434 1000 53502
rect 0 53378 94 53434
rect 150 53378 218 53434
rect 274 53378 342 53434
rect 398 53378 466 53434
rect 522 53378 590 53434
rect 646 53378 714 53434
rect 770 53378 838 53434
rect 894 53378 1000 53434
rect 0 53310 1000 53378
rect 0 53254 94 53310
rect 150 53254 218 53310
rect 274 53254 342 53310
rect 398 53254 466 53310
rect 522 53254 590 53310
rect 646 53254 714 53310
rect 770 53254 838 53310
rect 894 53254 1000 53310
rect 0 53186 1000 53254
rect 0 53130 94 53186
rect 150 53130 218 53186
rect 274 53130 342 53186
rect 398 53130 466 53186
rect 522 53130 590 53186
rect 646 53130 714 53186
rect 770 53130 838 53186
rect 894 53130 1000 53186
rect 0 53062 1000 53130
rect 0 53006 94 53062
rect 150 53006 218 53062
rect 274 53006 342 53062
rect 398 53006 466 53062
rect 522 53006 590 53062
rect 646 53006 714 53062
rect 770 53006 838 53062
rect 894 53006 1000 53062
rect 0 52938 1000 53006
rect 0 52882 94 52938
rect 150 52882 218 52938
rect 274 52882 342 52938
rect 398 52882 466 52938
rect 522 52882 590 52938
rect 646 52882 714 52938
rect 770 52882 838 52938
rect 894 52882 1000 52938
rect 0 52814 1000 52882
rect 0 52758 94 52814
rect 150 52758 218 52814
rect 274 52758 342 52814
rect 398 52758 466 52814
rect 522 52758 590 52814
rect 646 52758 714 52814
rect 770 52758 838 52814
rect 894 52758 1000 52814
rect 0 52690 1000 52758
rect 0 52634 94 52690
rect 150 52634 218 52690
rect 274 52634 342 52690
rect 398 52634 466 52690
rect 522 52634 590 52690
rect 646 52634 714 52690
rect 770 52634 838 52690
rect 894 52634 1000 52690
rect 0 52566 1000 52634
rect 0 52510 94 52566
rect 150 52510 218 52566
rect 274 52510 342 52566
rect 398 52510 466 52566
rect 522 52510 590 52566
rect 646 52510 714 52566
rect 770 52510 838 52566
rect 894 52510 1000 52566
rect 0 52400 1000 52510
rect 0 52079 1000 52200
rect 0 52023 94 52079
rect 150 52023 218 52079
rect 274 52023 342 52079
rect 398 52023 466 52079
rect 522 52023 590 52079
rect 646 52023 714 52079
rect 770 52023 838 52079
rect 894 52023 1000 52079
rect 0 51955 1000 52023
rect 0 51899 94 51955
rect 150 51899 218 51955
rect 274 51899 342 51955
rect 398 51899 466 51955
rect 522 51899 590 51955
rect 646 51899 714 51955
rect 770 51899 838 51955
rect 894 51899 1000 51955
rect 0 51831 1000 51899
rect 0 51775 94 51831
rect 150 51775 218 51831
rect 274 51775 342 51831
rect 398 51775 466 51831
rect 522 51775 590 51831
rect 646 51775 714 51831
rect 770 51775 838 51831
rect 894 51775 1000 51831
rect 0 51707 1000 51775
rect 0 51651 94 51707
rect 150 51651 218 51707
rect 274 51651 342 51707
rect 398 51651 466 51707
rect 522 51651 590 51707
rect 646 51651 714 51707
rect 770 51651 838 51707
rect 894 51651 1000 51707
rect 0 51583 1000 51651
rect 0 51527 94 51583
rect 150 51527 218 51583
rect 274 51527 342 51583
rect 398 51527 466 51583
rect 522 51527 590 51583
rect 646 51527 714 51583
rect 770 51527 838 51583
rect 894 51527 1000 51583
rect 0 51459 1000 51527
rect 0 51403 94 51459
rect 150 51403 218 51459
rect 274 51403 342 51459
rect 398 51403 466 51459
rect 522 51403 590 51459
rect 646 51403 714 51459
rect 770 51403 838 51459
rect 894 51403 1000 51459
rect 0 51335 1000 51403
rect 0 51279 94 51335
rect 150 51279 218 51335
rect 274 51279 342 51335
rect 398 51279 466 51335
rect 522 51279 590 51335
rect 646 51279 714 51335
rect 770 51279 838 51335
rect 894 51279 1000 51335
rect 0 51211 1000 51279
rect 0 51155 94 51211
rect 150 51155 218 51211
rect 274 51155 342 51211
rect 398 51155 466 51211
rect 522 51155 590 51211
rect 646 51155 714 51211
rect 770 51155 838 51211
rect 894 51155 1000 51211
rect 0 51087 1000 51155
rect 0 51031 94 51087
rect 150 51031 218 51087
rect 274 51031 342 51087
rect 398 51031 466 51087
rect 522 51031 590 51087
rect 646 51031 714 51087
rect 770 51031 838 51087
rect 894 51031 1000 51087
rect 0 50963 1000 51031
rect 0 50907 94 50963
rect 150 50907 218 50963
rect 274 50907 342 50963
rect 398 50907 466 50963
rect 522 50907 590 50963
rect 646 50907 714 50963
rect 770 50907 838 50963
rect 894 50907 1000 50963
rect 0 50800 1000 50907
rect 0 50480 1000 50600
rect 0 50424 95 50480
rect 151 50424 219 50480
rect 275 50424 343 50480
rect 399 50424 467 50480
rect 523 50424 591 50480
rect 647 50424 715 50480
rect 771 50424 839 50480
rect 895 50424 1000 50480
rect 0 50356 1000 50424
rect 0 50300 95 50356
rect 151 50300 219 50356
rect 275 50300 343 50356
rect 399 50300 467 50356
rect 523 50300 591 50356
rect 647 50300 715 50356
rect 771 50300 839 50356
rect 895 50300 1000 50356
rect 0 50232 1000 50300
rect 0 50176 95 50232
rect 151 50176 219 50232
rect 275 50176 343 50232
rect 399 50176 467 50232
rect 523 50176 591 50232
rect 647 50176 715 50232
rect 771 50176 839 50232
rect 895 50176 1000 50232
rect 0 50108 1000 50176
rect 0 50052 95 50108
rect 151 50052 219 50108
rect 275 50052 343 50108
rect 399 50052 467 50108
rect 523 50052 591 50108
rect 647 50052 715 50108
rect 771 50052 839 50108
rect 895 50052 1000 50108
rect 0 49984 1000 50052
rect 0 49928 95 49984
rect 151 49928 219 49984
rect 275 49928 343 49984
rect 399 49928 467 49984
rect 523 49928 591 49984
rect 647 49928 715 49984
rect 771 49928 839 49984
rect 895 49928 1000 49984
rect 0 49860 1000 49928
rect 0 49804 95 49860
rect 151 49804 219 49860
rect 275 49804 343 49860
rect 399 49804 467 49860
rect 523 49804 591 49860
rect 647 49804 715 49860
rect 771 49804 839 49860
rect 895 49804 1000 49860
rect 0 49736 1000 49804
rect 0 49680 95 49736
rect 151 49680 219 49736
rect 275 49680 343 49736
rect 399 49680 467 49736
rect 523 49680 591 49736
rect 647 49680 715 49736
rect 771 49680 839 49736
rect 895 49680 1000 49736
rect 0 49612 1000 49680
rect 0 49556 95 49612
rect 151 49556 219 49612
rect 275 49556 343 49612
rect 399 49556 467 49612
rect 523 49556 591 49612
rect 647 49556 715 49612
rect 771 49556 839 49612
rect 895 49556 1000 49612
rect 0 49488 1000 49556
rect 0 49432 95 49488
rect 151 49432 219 49488
rect 275 49432 343 49488
rect 399 49432 467 49488
rect 523 49432 591 49488
rect 647 49432 715 49488
rect 771 49432 839 49488
rect 895 49432 1000 49488
rect 0 49364 1000 49432
rect 0 49308 95 49364
rect 151 49308 219 49364
rect 275 49308 343 49364
rect 399 49308 467 49364
rect 523 49308 591 49364
rect 647 49308 715 49364
rect 771 49308 839 49364
rect 895 49308 1000 49364
rect 0 49200 1000 49308
rect 0 48893 1000 49000
rect 0 48837 94 48893
rect 150 48837 218 48893
rect 274 48837 342 48893
rect 398 48837 466 48893
rect 522 48837 590 48893
rect 646 48837 714 48893
rect 770 48837 838 48893
rect 894 48837 1000 48893
rect 0 48769 1000 48837
rect 0 48713 94 48769
rect 150 48713 218 48769
rect 274 48713 342 48769
rect 398 48713 466 48769
rect 522 48713 590 48769
rect 646 48713 714 48769
rect 770 48713 838 48769
rect 894 48713 1000 48769
rect 0 48645 1000 48713
rect 0 48589 94 48645
rect 150 48589 218 48645
rect 274 48589 342 48645
rect 398 48589 466 48645
rect 522 48589 590 48645
rect 646 48589 714 48645
rect 770 48589 838 48645
rect 894 48589 1000 48645
rect 0 48521 1000 48589
rect 0 48465 94 48521
rect 150 48465 218 48521
rect 274 48465 342 48521
rect 398 48465 466 48521
rect 522 48465 590 48521
rect 646 48465 714 48521
rect 770 48465 838 48521
rect 894 48465 1000 48521
rect 0 48397 1000 48465
rect 0 48341 94 48397
rect 150 48341 218 48397
rect 274 48341 342 48397
rect 398 48341 466 48397
rect 522 48341 590 48397
rect 646 48341 714 48397
rect 770 48341 838 48397
rect 894 48341 1000 48397
rect 0 48273 1000 48341
rect 0 48217 94 48273
rect 150 48217 218 48273
rect 274 48217 342 48273
rect 398 48217 466 48273
rect 522 48217 590 48273
rect 646 48217 714 48273
rect 770 48217 838 48273
rect 894 48217 1000 48273
rect 0 48149 1000 48217
rect 0 48093 94 48149
rect 150 48093 218 48149
rect 274 48093 342 48149
rect 398 48093 466 48149
rect 522 48093 590 48149
rect 646 48093 714 48149
rect 770 48093 838 48149
rect 894 48093 1000 48149
rect 0 48025 1000 48093
rect 0 47969 94 48025
rect 150 47969 218 48025
rect 274 47969 342 48025
rect 398 47969 466 48025
rect 522 47969 590 48025
rect 646 47969 714 48025
rect 770 47969 838 48025
rect 894 47969 1000 48025
rect 0 47901 1000 47969
rect 0 47845 94 47901
rect 150 47845 218 47901
rect 274 47845 342 47901
rect 398 47845 466 47901
rect 522 47845 590 47901
rect 646 47845 714 47901
rect 770 47845 838 47901
rect 894 47845 1000 47901
rect 0 47777 1000 47845
rect 0 47721 94 47777
rect 150 47721 218 47777
rect 274 47721 342 47777
rect 398 47721 466 47777
rect 522 47721 590 47777
rect 646 47721 714 47777
rect 770 47721 838 47777
rect 894 47721 1000 47777
rect 0 47653 1000 47721
rect 0 47597 94 47653
rect 150 47597 218 47653
rect 274 47597 342 47653
rect 398 47597 466 47653
rect 522 47597 590 47653
rect 646 47597 714 47653
rect 770 47597 838 47653
rect 894 47597 1000 47653
rect 0 47529 1000 47597
rect 0 47473 94 47529
rect 150 47473 218 47529
rect 274 47473 342 47529
rect 398 47473 466 47529
rect 522 47473 590 47529
rect 646 47473 714 47529
rect 770 47473 838 47529
rect 894 47473 1000 47529
rect 0 47405 1000 47473
rect 0 47349 94 47405
rect 150 47349 218 47405
rect 274 47349 342 47405
rect 398 47349 466 47405
rect 522 47349 590 47405
rect 646 47349 714 47405
rect 770 47349 838 47405
rect 894 47349 1000 47405
rect 0 47281 1000 47349
rect 0 47225 94 47281
rect 150 47225 218 47281
rect 274 47225 342 47281
rect 398 47225 466 47281
rect 522 47225 590 47281
rect 646 47225 714 47281
rect 770 47225 838 47281
rect 894 47225 1000 47281
rect 0 47157 1000 47225
rect 0 47101 94 47157
rect 150 47101 218 47157
rect 274 47101 342 47157
rect 398 47101 466 47157
rect 522 47101 590 47157
rect 646 47101 714 47157
rect 770 47101 838 47157
rect 894 47101 1000 47157
rect 0 47033 1000 47101
rect 0 46977 94 47033
rect 150 46977 218 47033
rect 274 46977 342 47033
rect 398 46977 466 47033
rect 522 46977 590 47033
rect 646 46977 714 47033
rect 770 46977 838 47033
rect 894 46977 1000 47033
rect 0 46909 1000 46977
rect 0 46853 94 46909
rect 150 46853 218 46909
rect 274 46853 342 46909
rect 398 46853 466 46909
rect 522 46853 590 46909
rect 646 46853 714 46909
rect 770 46853 838 46909
rect 894 46853 1000 46909
rect 0 46785 1000 46853
rect 0 46729 94 46785
rect 150 46729 218 46785
rect 274 46729 342 46785
rect 398 46729 466 46785
rect 522 46729 590 46785
rect 646 46729 714 46785
rect 770 46729 838 46785
rect 894 46729 1000 46785
rect 0 46661 1000 46729
rect 0 46605 94 46661
rect 150 46605 218 46661
rect 274 46605 342 46661
rect 398 46605 466 46661
rect 522 46605 590 46661
rect 646 46605 714 46661
rect 770 46605 838 46661
rect 894 46605 1000 46661
rect 0 46537 1000 46605
rect 0 46481 94 46537
rect 150 46481 218 46537
rect 274 46481 342 46537
rect 398 46481 466 46537
rect 522 46481 590 46537
rect 646 46481 714 46537
rect 770 46481 838 46537
rect 894 46481 1000 46537
rect 0 46413 1000 46481
rect 0 46357 94 46413
rect 150 46357 218 46413
rect 274 46357 342 46413
rect 398 46357 466 46413
rect 522 46357 590 46413
rect 646 46357 714 46413
rect 770 46357 838 46413
rect 894 46357 1000 46413
rect 0 46289 1000 46357
rect 0 46233 94 46289
rect 150 46233 218 46289
rect 274 46233 342 46289
rect 398 46233 466 46289
rect 522 46233 590 46289
rect 646 46233 714 46289
rect 770 46233 838 46289
rect 894 46233 1000 46289
rect 0 46165 1000 46233
rect 0 46109 94 46165
rect 150 46109 218 46165
rect 274 46109 342 46165
rect 398 46109 466 46165
rect 522 46109 590 46165
rect 646 46109 714 46165
rect 770 46109 838 46165
rect 894 46109 1000 46165
rect 0 46000 1000 46109
rect 0 45697 1000 45800
rect 0 45641 94 45697
rect 150 45641 218 45697
rect 274 45641 342 45697
rect 398 45641 466 45697
rect 522 45641 590 45697
rect 646 45641 714 45697
rect 770 45641 838 45697
rect 894 45641 1000 45697
rect 0 45573 1000 45641
rect 0 45517 94 45573
rect 150 45517 218 45573
rect 274 45517 342 45573
rect 398 45517 466 45573
rect 522 45517 590 45573
rect 646 45517 714 45573
rect 770 45517 838 45573
rect 894 45517 1000 45573
rect 0 45449 1000 45517
rect 0 45393 94 45449
rect 150 45393 218 45449
rect 274 45393 342 45449
rect 398 45393 466 45449
rect 522 45393 590 45449
rect 646 45393 714 45449
rect 770 45393 838 45449
rect 894 45393 1000 45449
rect 0 45325 1000 45393
rect 0 45269 94 45325
rect 150 45269 218 45325
rect 274 45269 342 45325
rect 398 45269 466 45325
rect 522 45269 590 45325
rect 646 45269 714 45325
rect 770 45269 838 45325
rect 894 45269 1000 45325
rect 0 45201 1000 45269
rect 0 45145 94 45201
rect 150 45145 218 45201
rect 274 45145 342 45201
rect 398 45145 466 45201
rect 522 45145 590 45201
rect 646 45145 714 45201
rect 770 45145 838 45201
rect 894 45145 1000 45201
rect 0 45077 1000 45145
rect 0 45021 94 45077
rect 150 45021 218 45077
rect 274 45021 342 45077
rect 398 45021 466 45077
rect 522 45021 590 45077
rect 646 45021 714 45077
rect 770 45021 838 45077
rect 894 45021 1000 45077
rect 0 44953 1000 45021
rect 0 44897 94 44953
rect 150 44897 218 44953
rect 274 44897 342 44953
rect 398 44897 466 44953
rect 522 44897 590 44953
rect 646 44897 714 44953
rect 770 44897 838 44953
rect 894 44897 1000 44953
rect 0 44829 1000 44897
rect 0 44773 94 44829
rect 150 44773 218 44829
rect 274 44773 342 44829
rect 398 44773 466 44829
rect 522 44773 590 44829
rect 646 44773 714 44829
rect 770 44773 838 44829
rect 894 44773 1000 44829
rect 0 44705 1000 44773
rect 0 44649 94 44705
rect 150 44649 218 44705
rect 274 44649 342 44705
rect 398 44649 466 44705
rect 522 44649 590 44705
rect 646 44649 714 44705
rect 770 44649 838 44705
rect 894 44649 1000 44705
rect 0 44581 1000 44649
rect 0 44525 94 44581
rect 150 44525 218 44581
rect 274 44525 342 44581
rect 398 44525 466 44581
rect 522 44525 590 44581
rect 646 44525 714 44581
rect 770 44525 838 44581
rect 894 44525 1000 44581
rect 0 44457 1000 44525
rect 0 44401 94 44457
rect 150 44401 218 44457
rect 274 44401 342 44457
rect 398 44401 466 44457
rect 522 44401 590 44457
rect 646 44401 714 44457
rect 770 44401 838 44457
rect 894 44401 1000 44457
rect 0 44333 1000 44401
rect 0 44277 94 44333
rect 150 44277 218 44333
rect 274 44277 342 44333
rect 398 44277 466 44333
rect 522 44277 590 44333
rect 646 44277 714 44333
rect 770 44277 838 44333
rect 894 44277 1000 44333
rect 0 44209 1000 44277
rect 0 44153 94 44209
rect 150 44153 218 44209
rect 274 44153 342 44209
rect 398 44153 466 44209
rect 522 44153 590 44209
rect 646 44153 714 44209
rect 770 44153 838 44209
rect 894 44153 1000 44209
rect 0 44085 1000 44153
rect 0 44029 94 44085
rect 150 44029 218 44085
rect 274 44029 342 44085
rect 398 44029 466 44085
rect 522 44029 590 44085
rect 646 44029 714 44085
rect 770 44029 838 44085
rect 894 44029 1000 44085
rect 0 43961 1000 44029
rect 0 43905 94 43961
rect 150 43905 218 43961
rect 274 43905 342 43961
rect 398 43905 466 43961
rect 522 43905 590 43961
rect 646 43905 714 43961
rect 770 43905 838 43961
rect 894 43905 1000 43961
rect 0 43837 1000 43905
rect 0 43781 94 43837
rect 150 43781 218 43837
rect 274 43781 342 43837
rect 398 43781 466 43837
rect 522 43781 590 43837
rect 646 43781 714 43837
rect 770 43781 838 43837
rect 894 43781 1000 43837
rect 0 43713 1000 43781
rect 0 43657 94 43713
rect 150 43657 218 43713
rect 274 43657 342 43713
rect 398 43657 466 43713
rect 522 43657 590 43713
rect 646 43657 714 43713
rect 770 43657 838 43713
rect 894 43657 1000 43713
rect 0 43589 1000 43657
rect 0 43533 94 43589
rect 150 43533 218 43589
rect 274 43533 342 43589
rect 398 43533 466 43589
rect 522 43533 590 43589
rect 646 43533 714 43589
rect 770 43533 838 43589
rect 894 43533 1000 43589
rect 0 43465 1000 43533
rect 0 43409 94 43465
rect 150 43409 218 43465
rect 274 43409 342 43465
rect 398 43409 466 43465
rect 522 43409 590 43465
rect 646 43409 714 43465
rect 770 43409 838 43465
rect 894 43409 1000 43465
rect 0 43341 1000 43409
rect 0 43285 94 43341
rect 150 43285 218 43341
rect 274 43285 342 43341
rect 398 43285 466 43341
rect 522 43285 590 43341
rect 646 43285 714 43341
rect 770 43285 838 43341
rect 894 43285 1000 43341
rect 0 43217 1000 43285
rect 0 43161 94 43217
rect 150 43161 218 43217
rect 274 43161 342 43217
rect 398 43161 466 43217
rect 522 43161 590 43217
rect 646 43161 714 43217
rect 770 43161 838 43217
rect 894 43161 1000 43217
rect 0 43093 1000 43161
rect 0 43037 94 43093
rect 150 43037 218 43093
rect 274 43037 342 43093
rect 398 43037 466 43093
rect 522 43037 590 43093
rect 646 43037 714 43093
rect 770 43037 838 43093
rect 894 43037 1000 43093
rect 0 42969 1000 43037
rect 0 42913 94 42969
rect 150 42913 218 42969
rect 274 42913 342 42969
rect 398 42913 466 42969
rect 522 42913 590 42969
rect 646 42913 714 42969
rect 770 42913 838 42969
rect 894 42913 1000 42969
rect 0 42800 1000 42913
rect 0 42484 1000 42600
rect 0 42428 95 42484
rect 151 42428 219 42484
rect 275 42428 343 42484
rect 399 42428 467 42484
rect 523 42428 591 42484
rect 647 42428 715 42484
rect 771 42428 839 42484
rect 895 42428 1000 42484
rect 0 42360 1000 42428
rect 0 42304 95 42360
rect 151 42304 219 42360
rect 275 42304 343 42360
rect 399 42304 467 42360
rect 523 42304 591 42360
rect 647 42304 715 42360
rect 771 42304 839 42360
rect 895 42304 1000 42360
rect 0 42236 1000 42304
rect 0 42180 95 42236
rect 151 42180 219 42236
rect 275 42180 343 42236
rect 399 42180 467 42236
rect 523 42180 591 42236
rect 647 42180 715 42236
rect 771 42180 839 42236
rect 895 42180 1000 42236
rect 0 42112 1000 42180
rect 0 42056 95 42112
rect 151 42056 219 42112
rect 275 42056 343 42112
rect 399 42056 467 42112
rect 523 42056 591 42112
rect 647 42056 715 42112
rect 771 42056 839 42112
rect 895 42056 1000 42112
rect 0 41988 1000 42056
rect 0 41932 95 41988
rect 151 41932 219 41988
rect 275 41932 343 41988
rect 399 41932 467 41988
rect 523 41932 591 41988
rect 647 41932 715 41988
rect 771 41932 839 41988
rect 895 41932 1000 41988
rect 0 41864 1000 41932
rect 0 41808 95 41864
rect 151 41808 219 41864
rect 275 41808 343 41864
rect 399 41808 467 41864
rect 523 41808 591 41864
rect 647 41808 715 41864
rect 771 41808 839 41864
rect 895 41808 1000 41864
rect 0 41740 1000 41808
rect 0 41684 95 41740
rect 151 41684 219 41740
rect 275 41684 343 41740
rect 399 41684 467 41740
rect 523 41684 591 41740
rect 647 41684 715 41740
rect 771 41684 839 41740
rect 895 41684 1000 41740
rect 0 41616 1000 41684
rect 0 41560 95 41616
rect 151 41560 219 41616
rect 275 41560 343 41616
rect 399 41560 467 41616
rect 523 41560 591 41616
rect 647 41560 715 41616
rect 771 41560 839 41616
rect 895 41560 1000 41616
rect 0 41492 1000 41560
rect 0 41436 95 41492
rect 151 41436 219 41492
rect 275 41436 343 41492
rect 399 41436 467 41492
rect 523 41436 591 41492
rect 647 41436 715 41492
rect 771 41436 839 41492
rect 895 41436 1000 41492
rect 0 41368 1000 41436
rect 0 41312 95 41368
rect 151 41312 219 41368
rect 275 41312 343 41368
rect 399 41312 467 41368
rect 523 41312 591 41368
rect 647 41312 715 41368
rect 771 41312 839 41368
rect 895 41312 1000 41368
rect 0 41200 1000 41312
rect 0 40896 1000 41000
rect 0 40840 95 40896
rect 151 40840 219 40896
rect 275 40840 343 40896
rect 399 40840 467 40896
rect 523 40840 591 40896
rect 647 40840 715 40896
rect 771 40840 839 40896
rect 895 40840 1000 40896
rect 0 40772 1000 40840
rect 0 40716 95 40772
rect 151 40716 219 40772
rect 275 40716 343 40772
rect 399 40716 467 40772
rect 523 40716 591 40772
rect 647 40716 715 40772
rect 771 40716 839 40772
rect 895 40716 1000 40772
rect 0 40648 1000 40716
rect 0 40592 95 40648
rect 151 40592 219 40648
rect 275 40592 343 40648
rect 399 40592 467 40648
rect 523 40592 591 40648
rect 647 40592 715 40648
rect 771 40592 839 40648
rect 895 40592 1000 40648
rect 0 40524 1000 40592
rect 0 40468 95 40524
rect 151 40468 219 40524
rect 275 40468 343 40524
rect 399 40468 467 40524
rect 523 40468 591 40524
rect 647 40468 715 40524
rect 771 40468 839 40524
rect 895 40468 1000 40524
rect 0 40400 1000 40468
rect 0 40344 95 40400
rect 151 40344 219 40400
rect 275 40344 343 40400
rect 399 40344 467 40400
rect 523 40344 591 40400
rect 647 40344 715 40400
rect 771 40344 839 40400
rect 895 40344 1000 40400
rect 0 40276 1000 40344
rect 0 40220 95 40276
rect 151 40220 219 40276
rect 275 40220 343 40276
rect 399 40220 467 40276
rect 523 40220 591 40276
rect 647 40220 715 40276
rect 771 40220 839 40276
rect 895 40220 1000 40276
rect 0 40152 1000 40220
rect 0 40096 95 40152
rect 151 40096 219 40152
rect 275 40096 343 40152
rect 399 40096 467 40152
rect 523 40096 591 40152
rect 647 40096 715 40152
rect 771 40096 839 40152
rect 895 40096 1000 40152
rect 0 40028 1000 40096
rect 0 39972 95 40028
rect 151 39972 219 40028
rect 275 39972 343 40028
rect 399 39972 467 40028
rect 523 39972 591 40028
rect 647 39972 715 40028
rect 771 39972 839 40028
rect 895 39972 1000 40028
rect 0 39904 1000 39972
rect 0 39848 95 39904
rect 151 39848 219 39904
rect 275 39848 343 39904
rect 399 39848 467 39904
rect 523 39848 591 39904
rect 647 39848 715 39904
rect 771 39848 839 39904
rect 895 39848 1000 39904
rect 0 39780 1000 39848
rect 0 39724 95 39780
rect 151 39724 219 39780
rect 275 39724 343 39780
rect 399 39724 467 39780
rect 523 39724 591 39780
rect 647 39724 715 39780
rect 771 39724 839 39780
rect 895 39724 1000 39780
rect 0 39600 1000 39724
rect 0 39304 1000 39400
rect 0 39248 94 39304
rect 150 39248 218 39304
rect 274 39248 342 39304
rect 398 39248 466 39304
rect 522 39248 590 39304
rect 646 39248 714 39304
rect 770 39248 838 39304
rect 894 39248 1000 39304
rect 0 39180 1000 39248
rect 0 39124 94 39180
rect 150 39124 218 39180
rect 274 39124 342 39180
rect 398 39124 466 39180
rect 522 39124 590 39180
rect 646 39124 714 39180
rect 770 39124 838 39180
rect 894 39124 1000 39180
rect 0 39056 1000 39124
rect 0 39000 94 39056
rect 150 39000 218 39056
rect 274 39000 342 39056
rect 398 39000 466 39056
rect 522 39000 590 39056
rect 646 39000 714 39056
rect 770 39000 838 39056
rect 894 39000 1000 39056
rect 0 38932 1000 39000
rect 0 38876 94 38932
rect 150 38876 218 38932
rect 274 38876 342 38932
rect 398 38876 466 38932
rect 522 38876 590 38932
rect 646 38876 714 38932
rect 770 38876 838 38932
rect 894 38876 1000 38932
rect 0 38808 1000 38876
rect 0 38752 94 38808
rect 150 38752 218 38808
rect 274 38752 342 38808
rect 398 38752 466 38808
rect 522 38752 590 38808
rect 646 38752 714 38808
rect 770 38752 838 38808
rect 894 38752 1000 38808
rect 0 38684 1000 38752
rect 0 38628 94 38684
rect 150 38628 218 38684
rect 274 38628 342 38684
rect 398 38628 466 38684
rect 522 38628 590 38684
rect 646 38628 714 38684
rect 770 38628 838 38684
rect 894 38628 1000 38684
rect 0 38560 1000 38628
rect 0 38504 94 38560
rect 150 38504 218 38560
rect 274 38504 342 38560
rect 398 38504 466 38560
rect 522 38504 590 38560
rect 646 38504 714 38560
rect 770 38504 838 38560
rect 894 38504 1000 38560
rect 0 38436 1000 38504
rect 0 38380 94 38436
rect 150 38380 218 38436
rect 274 38380 342 38436
rect 398 38380 466 38436
rect 522 38380 590 38436
rect 646 38380 714 38436
rect 770 38380 838 38436
rect 894 38380 1000 38436
rect 0 38312 1000 38380
rect 0 38256 94 38312
rect 150 38256 218 38312
rect 274 38256 342 38312
rect 398 38256 466 38312
rect 522 38256 590 38312
rect 646 38256 714 38312
rect 770 38256 838 38312
rect 894 38256 1000 38312
rect 0 38188 1000 38256
rect 0 38132 94 38188
rect 150 38132 218 38188
rect 274 38132 342 38188
rect 398 38132 466 38188
rect 522 38132 590 38188
rect 646 38132 714 38188
rect 770 38132 838 38188
rect 894 38132 1000 38188
rect 0 38064 1000 38132
rect 0 38008 94 38064
rect 150 38008 218 38064
rect 274 38008 342 38064
rect 398 38008 466 38064
rect 522 38008 590 38064
rect 646 38008 714 38064
rect 770 38008 838 38064
rect 894 38008 1000 38064
rect 0 37940 1000 38008
rect 0 37884 94 37940
rect 150 37884 218 37940
rect 274 37884 342 37940
rect 398 37884 466 37940
rect 522 37884 590 37940
rect 646 37884 714 37940
rect 770 37884 838 37940
rect 894 37884 1000 37940
rect 0 37816 1000 37884
rect 0 37760 94 37816
rect 150 37760 218 37816
rect 274 37760 342 37816
rect 398 37760 466 37816
rect 522 37760 590 37816
rect 646 37760 714 37816
rect 770 37760 838 37816
rect 894 37760 1000 37816
rect 0 37692 1000 37760
rect 0 37636 94 37692
rect 150 37636 218 37692
rect 274 37636 342 37692
rect 398 37636 466 37692
rect 522 37636 590 37692
rect 646 37636 714 37692
rect 770 37636 838 37692
rect 894 37636 1000 37692
rect 0 37568 1000 37636
rect 0 37512 94 37568
rect 150 37512 218 37568
rect 274 37512 342 37568
rect 398 37512 466 37568
rect 522 37512 590 37568
rect 646 37512 714 37568
rect 770 37512 838 37568
rect 894 37512 1000 37568
rect 0 37444 1000 37512
rect 0 37388 94 37444
rect 150 37388 218 37444
rect 274 37388 342 37444
rect 398 37388 466 37444
rect 522 37388 590 37444
rect 646 37388 714 37444
rect 770 37388 838 37444
rect 894 37388 1000 37444
rect 0 37320 1000 37388
rect 0 37264 94 37320
rect 150 37264 218 37320
rect 274 37264 342 37320
rect 398 37264 466 37320
rect 522 37264 590 37320
rect 646 37264 714 37320
rect 770 37264 838 37320
rect 894 37264 1000 37320
rect 0 37196 1000 37264
rect 0 37140 94 37196
rect 150 37140 218 37196
rect 274 37140 342 37196
rect 398 37140 466 37196
rect 522 37140 590 37196
rect 646 37140 714 37196
rect 770 37140 838 37196
rect 894 37140 1000 37196
rect 0 37072 1000 37140
rect 0 37016 94 37072
rect 150 37016 218 37072
rect 274 37016 342 37072
rect 398 37016 466 37072
rect 522 37016 590 37072
rect 646 37016 714 37072
rect 770 37016 838 37072
rect 894 37016 1000 37072
rect 0 36948 1000 37016
rect 0 36892 94 36948
rect 150 36892 218 36948
rect 274 36892 342 36948
rect 398 36892 466 36948
rect 522 36892 590 36948
rect 646 36892 714 36948
rect 770 36892 838 36948
rect 894 36892 1000 36948
rect 0 36824 1000 36892
rect 0 36768 94 36824
rect 150 36768 218 36824
rect 274 36768 342 36824
rect 398 36768 466 36824
rect 522 36768 590 36824
rect 646 36768 714 36824
rect 770 36768 838 36824
rect 894 36768 1000 36824
rect 0 36700 1000 36768
rect 0 36644 94 36700
rect 150 36644 218 36700
rect 274 36644 342 36700
rect 398 36644 466 36700
rect 522 36644 590 36700
rect 646 36644 714 36700
rect 770 36644 838 36700
rect 894 36644 1000 36700
rect 0 36576 1000 36644
rect 0 36520 94 36576
rect 150 36520 218 36576
rect 274 36520 342 36576
rect 398 36520 466 36576
rect 522 36520 590 36576
rect 646 36520 714 36576
rect 770 36520 838 36576
rect 894 36520 1000 36576
rect 0 36400 1000 36520
rect 0 36094 1000 36200
rect 0 36038 94 36094
rect 150 36038 218 36094
rect 274 36038 342 36094
rect 398 36038 466 36094
rect 522 36038 590 36094
rect 646 36038 714 36094
rect 770 36038 838 36094
rect 894 36038 1000 36094
rect 0 35970 1000 36038
rect 0 35914 94 35970
rect 150 35914 218 35970
rect 274 35914 342 35970
rect 398 35914 466 35970
rect 522 35914 590 35970
rect 646 35914 714 35970
rect 770 35914 838 35970
rect 894 35914 1000 35970
rect 0 35846 1000 35914
rect 0 35790 94 35846
rect 150 35790 218 35846
rect 274 35790 342 35846
rect 398 35790 466 35846
rect 522 35790 590 35846
rect 646 35790 714 35846
rect 770 35790 838 35846
rect 894 35790 1000 35846
rect 0 35722 1000 35790
rect 0 35666 94 35722
rect 150 35666 218 35722
rect 274 35666 342 35722
rect 398 35666 466 35722
rect 522 35666 590 35722
rect 646 35666 714 35722
rect 770 35666 838 35722
rect 894 35666 1000 35722
rect 0 35598 1000 35666
rect 0 35542 94 35598
rect 150 35542 218 35598
rect 274 35542 342 35598
rect 398 35542 466 35598
rect 522 35542 590 35598
rect 646 35542 714 35598
rect 770 35542 838 35598
rect 894 35542 1000 35598
rect 0 35474 1000 35542
rect 0 35418 94 35474
rect 150 35418 218 35474
rect 274 35418 342 35474
rect 398 35418 466 35474
rect 522 35418 590 35474
rect 646 35418 714 35474
rect 770 35418 838 35474
rect 894 35418 1000 35474
rect 0 35350 1000 35418
rect 0 35294 94 35350
rect 150 35294 218 35350
rect 274 35294 342 35350
rect 398 35294 466 35350
rect 522 35294 590 35350
rect 646 35294 714 35350
rect 770 35294 838 35350
rect 894 35294 1000 35350
rect 0 35226 1000 35294
rect 0 35170 94 35226
rect 150 35170 218 35226
rect 274 35170 342 35226
rect 398 35170 466 35226
rect 522 35170 590 35226
rect 646 35170 714 35226
rect 770 35170 838 35226
rect 894 35170 1000 35226
rect 0 35102 1000 35170
rect 0 35046 94 35102
rect 150 35046 218 35102
rect 274 35046 342 35102
rect 398 35046 466 35102
rect 522 35046 590 35102
rect 646 35046 714 35102
rect 770 35046 838 35102
rect 894 35046 1000 35102
rect 0 34978 1000 35046
rect 0 34922 94 34978
rect 150 34922 218 34978
rect 274 34922 342 34978
rect 398 34922 466 34978
rect 522 34922 590 34978
rect 646 34922 714 34978
rect 770 34922 838 34978
rect 894 34922 1000 34978
rect 0 34854 1000 34922
rect 0 34798 94 34854
rect 150 34798 218 34854
rect 274 34798 342 34854
rect 398 34798 466 34854
rect 522 34798 590 34854
rect 646 34798 714 34854
rect 770 34798 838 34854
rect 894 34798 1000 34854
rect 0 34730 1000 34798
rect 0 34674 94 34730
rect 150 34674 218 34730
rect 274 34674 342 34730
rect 398 34674 466 34730
rect 522 34674 590 34730
rect 646 34674 714 34730
rect 770 34674 838 34730
rect 894 34674 1000 34730
rect 0 34606 1000 34674
rect 0 34550 94 34606
rect 150 34550 218 34606
rect 274 34550 342 34606
rect 398 34550 466 34606
rect 522 34550 590 34606
rect 646 34550 714 34606
rect 770 34550 838 34606
rect 894 34550 1000 34606
rect 0 34482 1000 34550
rect 0 34426 94 34482
rect 150 34426 218 34482
rect 274 34426 342 34482
rect 398 34426 466 34482
rect 522 34426 590 34482
rect 646 34426 714 34482
rect 770 34426 838 34482
rect 894 34426 1000 34482
rect 0 34358 1000 34426
rect 0 34302 94 34358
rect 150 34302 218 34358
rect 274 34302 342 34358
rect 398 34302 466 34358
rect 522 34302 590 34358
rect 646 34302 714 34358
rect 770 34302 838 34358
rect 894 34302 1000 34358
rect 0 34234 1000 34302
rect 0 34178 94 34234
rect 150 34178 218 34234
rect 274 34178 342 34234
rect 398 34178 466 34234
rect 522 34178 590 34234
rect 646 34178 714 34234
rect 770 34178 838 34234
rect 894 34178 1000 34234
rect 0 34110 1000 34178
rect 0 34054 94 34110
rect 150 34054 218 34110
rect 274 34054 342 34110
rect 398 34054 466 34110
rect 522 34054 590 34110
rect 646 34054 714 34110
rect 770 34054 838 34110
rect 894 34054 1000 34110
rect 0 33986 1000 34054
rect 0 33930 94 33986
rect 150 33930 218 33986
rect 274 33930 342 33986
rect 398 33930 466 33986
rect 522 33930 590 33986
rect 646 33930 714 33986
rect 770 33930 838 33986
rect 894 33930 1000 33986
rect 0 33862 1000 33930
rect 0 33806 94 33862
rect 150 33806 218 33862
rect 274 33806 342 33862
rect 398 33806 466 33862
rect 522 33806 590 33862
rect 646 33806 714 33862
rect 770 33806 838 33862
rect 894 33806 1000 33862
rect 0 33738 1000 33806
rect 0 33682 94 33738
rect 150 33682 218 33738
rect 274 33682 342 33738
rect 398 33682 466 33738
rect 522 33682 590 33738
rect 646 33682 714 33738
rect 770 33682 838 33738
rect 894 33682 1000 33738
rect 0 33614 1000 33682
rect 0 33558 94 33614
rect 150 33558 218 33614
rect 274 33558 342 33614
rect 398 33558 466 33614
rect 522 33558 590 33614
rect 646 33558 714 33614
rect 770 33558 838 33614
rect 894 33558 1000 33614
rect 0 33490 1000 33558
rect 0 33434 94 33490
rect 150 33434 218 33490
rect 274 33434 342 33490
rect 398 33434 466 33490
rect 522 33434 590 33490
rect 646 33434 714 33490
rect 770 33434 838 33490
rect 894 33434 1000 33490
rect 0 33366 1000 33434
rect 0 33310 94 33366
rect 150 33310 218 33366
rect 274 33310 342 33366
rect 398 33310 466 33366
rect 522 33310 590 33366
rect 646 33310 714 33366
rect 770 33310 838 33366
rect 894 33310 1000 33366
rect 0 33200 1000 33310
rect 0 32902 1000 33000
rect 0 32846 94 32902
rect 150 32846 218 32902
rect 274 32846 342 32902
rect 398 32846 466 32902
rect 522 32846 590 32902
rect 646 32846 714 32902
rect 770 32846 838 32902
rect 894 32846 1000 32902
rect 0 32778 1000 32846
rect 0 32722 94 32778
rect 150 32722 218 32778
rect 274 32722 342 32778
rect 398 32722 466 32778
rect 522 32722 590 32778
rect 646 32722 714 32778
rect 770 32722 838 32778
rect 894 32722 1000 32778
rect 0 32654 1000 32722
rect 0 32598 94 32654
rect 150 32598 218 32654
rect 274 32598 342 32654
rect 398 32598 466 32654
rect 522 32598 590 32654
rect 646 32598 714 32654
rect 770 32598 838 32654
rect 894 32598 1000 32654
rect 0 32530 1000 32598
rect 0 32474 94 32530
rect 150 32474 218 32530
rect 274 32474 342 32530
rect 398 32474 466 32530
rect 522 32474 590 32530
rect 646 32474 714 32530
rect 770 32474 838 32530
rect 894 32474 1000 32530
rect 0 32406 1000 32474
rect 0 32350 94 32406
rect 150 32350 218 32406
rect 274 32350 342 32406
rect 398 32350 466 32406
rect 522 32350 590 32406
rect 646 32350 714 32406
rect 770 32350 838 32406
rect 894 32350 1000 32406
rect 0 32282 1000 32350
rect 0 32226 94 32282
rect 150 32226 218 32282
rect 274 32226 342 32282
rect 398 32226 466 32282
rect 522 32226 590 32282
rect 646 32226 714 32282
rect 770 32226 838 32282
rect 894 32226 1000 32282
rect 0 32158 1000 32226
rect 0 32102 94 32158
rect 150 32102 218 32158
rect 274 32102 342 32158
rect 398 32102 466 32158
rect 522 32102 590 32158
rect 646 32102 714 32158
rect 770 32102 838 32158
rect 894 32102 1000 32158
rect 0 32034 1000 32102
rect 0 31978 94 32034
rect 150 31978 218 32034
rect 274 31978 342 32034
rect 398 31978 466 32034
rect 522 31978 590 32034
rect 646 31978 714 32034
rect 770 31978 838 32034
rect 894 31978 1000 32034
rect 0 31910 1000 31978
rect 0 31854 94 31910
rect 150 31854 218 31910
rect 274 31854 342 31910
rect 398 31854 466 31910
rect 522 31854 590 31910
rect 646 31854 714 31910
rect 770 31854 838 31910
rect 894 31854 1000 31910
rect 0 31786 1000 31854
rect 0 31730 94 31786
rect 150 31730 218 31786
rect 274 31730 342 31786
rect 398 31730 466 31786
rect 522 31730 590 31786
rect 646 31730 714 31786
rect 770 31730 838 31786
rect 894 31730 1000 31786
rect 0 31662 1000 31730
rect 0 31606 94 31662
rect 150 31606 218 31662
rect 274 31606 342 31662
rect 398 31606 466 31662
rect 522 31606 590 31662
rect 646 31606 714 31662
rect 770 31606 838 31662
rect 894 31606 1000 31662
rect 0 31538 1000 31606
rect 0 31482 94 31538
rect 150 31482 218 31538
rect 274 31482 342 31538
rect 398 31482 466 31538
rect 522 31482 590 31538
rect 646 31482 714 31538
rect 770 31482 838 31538
rect 894 31482 1000 31538
rect 0 31414 1000 31482
rect 0 31358 94 31414
rect 150 31358 218 31414
rect 274 31358 342 31414
rect 398 31358 466 31414
rect 522 31358 590 31414
rect 646 31358 714 31414
rect 770 31358 838 31414
rect 894 31358 1000 31414
rect 0 31290 1000 31358
rect 0 31234 94 31290
rect 150 31234 218 31290
rect 274 31234 342 31290
rect 398 31234 466 31290
rect 522 31234 590 31290
rect 646 31234 714 31290
rect 770 31234 838 31290
rect 894 31234 1000 31290
rect 0 31166 1000 31234
rect 0 31110 94 31166
rect 150 31110 218 31166
rect 274 31110 342 31166
rect 398 31110 466 31166
rect 522 31110 590 31166
rect 646 31110 714 31166
rect 770 31110 838 31166
rect 894 31110 1000 31166
rect 0 31042 1000 31110
rect 0 30986 94 31042
rect 150 30986 218 31042
rect 274 30986 342 31042
rect 398 30986 466 31042
rect 522 30986 590 31042
rect 646 30986 714 31042
rect 770 30986 838 31042
rect 894 30986 1000 31042
rect 0 30918 1000 30986
rect 0 30862 94 30918
rect 150 30862 218 30918
rect 274 30862 342 30918
rect 398 30862 466 30918
rect 522 30862 590 30918
rect 646 30862 714 30918
rect 770 30862 838 30918
rect 894 30862 1000 30918
rect 0 30794 1000 30862
rect 0 30738 94 30794
rect 150 30738 218 30794
rect 274 30738 342 30794
rect 398 30738 466 30794
rect 522 30738 590 30794
rect 646 30738 714 30794
rect 770 30738 838 30794
rect 894 30738 1000 30794
rect 0 30670 1000 30738
rect 0 30614 94 30670
rect 150 30614 218 30670
rect 274 30614 342 30670
rect 398 30614 466 30670
rect 522 30614 590 30670
rect 646 30614 714 30670
rect 770 30614 838 30670
rect 894 30614 1000 30670
rect 0 30546 1000 30614
rect 0 30490 94 30546
rect 150 30490 218 30546
rect 274 30490 342 30546
rect 398 30490 466 30546
rect 522 30490 590 30546
rect 646 30490 714 30546
rect 770 30490 838 30546
rect 894 30490 1000 30546
rect 0 30422 1000 30490
rect 0 30366 94 30422
rect 150 30366 218 30422
rect 274 30366 342 30422
rect 398 30366 466 30422
rect 522 30366 590 30422
rect 646 30366 714 30422
rect 770 30366 838 30422
rect 894 30366 1000 30422
rect 0 30298 1000 30366
rect 0 30242 94 30298
rect 150 30242 218 30298
rect 274 30242 342 30298
rect 398 30242 466 30298
rect 522 30242 590 30298
rect 646 30242 714 30298
rect 770 30242 838 30298
rect 894 30242 1000 30298
rect 0 30174 1000 30242
rect 0 30118 94 30174
rect 150 30118 218 30174
rect 274 30118 342 30174
rect 398 30118 466 30174
rect 522 30118 590 30174
rect 646 30118 714 30174
rect 770 30118 838 30174
rect 894 30118 1000 30174
rect 0 30000 1000 30118
rect 0 29685 1000 29800
rect 0 29629 94 29685
rect 150 29629 218 29685
rect 274 29629 342 29685
rect 398 29629 466 29685
rect 522 29629 590 29685
rect 646 29629 714 29685
rect 770 29629 838 29685
rect 894 29629 1000 29685
rect 0 29561 1000 29629
rect 0 29505 94 29561
rect 150 29505 218 29561
rect 274 29505 342 29561
rect 398 29505 466 29561
rect 522 29505 590 29561
rect 646 29505 714 29561
rect 770 29505 838 29561
rect 894 29505 1000 29561
rect 0 29437 1000 29505
rect 0 29381 94 29437
rect 150 29381 218 29437
rect 274 29381 342 29437
rect 398 29381 466 29437
rect 522 29381 590 29437
rect 646 29381 714 29437
rect 770 29381 838 29437
rect 894 29381 1000 29437
rect 0 29313 1000 29381
rect 0 29257 94 29313
rect 150 29257 218 29313
rect 274 29257 342 29313
rect 398 29257 466 29313
rect 522 29257 590 29313
rect 646 29257 714 29313
rect 770 29257 838 29313
rect 894 29257 1000 29313
rect 0 29189 1000 29257
rect 0 29133 94 29189
rect 150 29133 218 29189
rect 274 29133 342 29189
rect 398 29133 466 29189
rect 522 29133 590 29189
rect 646 29133 714 29189
rect 770 29133 838 29189
rect 894 29133 1000 29189
rect 0 29065 1000 29133
rect 0 29009 94 29065
rect 150 29009 218 29065
rect 274 29009 342 29065
rect 398 29009 466 29065
rect 522 29009 590 29065
rect 646 29009 714 29065
rect 770 29009 838 29065
rect 894 29009 1000 29065
rect 0 28941 1000 29009
rect 0 28885 94 28941
rect 150 28885 218 28941
rect 274 28885 342 28941
rect 398 28885 466 28941
rect 522 28885 590 28941
rect 646 28885 714 28941
rect 770 28885 838 28941
rect 894 28885 1000 28941
rect 0 28817 1000 28885
rect 0 28761 94 28817
rect 150 28761 218 28817
rect 274 28761 342 28817
rect 398 28761 466 28817
rect 522 28761 590 28817
rect 646 28761 714 28817
rect 770 28761 838 28817
rect 894 28761 1000 28817
rect 0 28693 1000 28761
rect 0 28637 94 28693
rect 150 28637 218 28693
rect 274 28637 342 28693
rect 398 28637 466 28693
rect 522 28637 590 28693
rect 646 28637 714 28693
rect 770 28637 838 28693
rect 894 28637 1000 28693
rect 0 28569 1000 28637
rect 0 28513 94 28569
rect 150 28513 218 28569
rect 274 28513 342 28569
rect 398 28513 466 28569
rect 522 28513 590 28569
rect 646 28513 714 28569
rect 770 28513 838 28569
rect 894 28513 1000 28569
rect 0 28445 1000 28513
rect 0 28389 94 28445
rect 150 28389 218 28445
rect 274 28389 342 28445
rect 398 28389 466 28445
rect 522 28389 590 28445
rect 646 28389 714 28445
rect 770 28389 838 28445
rect 894 28389 1000 28445
rect 0 28321 1000 28389
rect 0 28265 94 28321
rect 150 28265 218 28321
rect 274 28265 342 28321
rect 398 28265 466 28321
rect 522 28265 590 28321
rect 646 28265 714 28321
rect 770 28265 838 28321
rect 894 28265 1000 28321
rect 0 28197 1000 28265
rect 0 28141 94 28197
rect 150 28141 218 28197
rect 274 28141 342 28197
rect 398 28141 466 28197
rect 522 28141 590 28197
rect 646 28141 714 28197
rect 770 28141 838 28197
rect 894 28141 1000 28197
rect 0 28073 1000 28141
rect 0 28017 94 28073
rect 150 28017 218 28073
rect 274 28017 342 28073
rect 398 28017 466 28073
rect 522 28017 590 28073
rect 646 28017 714 28073
rect 770 28017 838 28073
rect 894 28017 1000 28073
rect 0 27949 1000 28017
rect 0 27893 94 27949
rect 150 27893 218 27949
rect 274 27893 342 27949
rect 398 27893 466 27949
rect 522 27893 590 27949
rect 646 27893 714 27949
rect 770 27893 838 27949
rect 894 27893 1000 27949
rect 0 27825 1000 27893
rect 0 27769 94 27825
rect 150 27769 218 27825
rect 274 27769 342 27825
rect 398 27769 466 27825
rect 522 27769 590 27825
rect 646 27769 714 27825
rect 770 27769 838 27825
rect 894 27769 1000 27825
rect 0 27701 1000 27769
rect 0 27645 94 27701
rect 150 27645 218 27701
rect 274 27645 342 27701
rect 398 27645 466 27701
rect 522 27645 590 27701
rect 646 27645 714 27701
rect 770 27645 838 27701
rect 894 27645 1000 27701
rect 0 27577 1000 27645
rect 0 27521 94 27577
rect 150 27521 218 27577
rect 274 27521 342 27577
rect 398 27521 466 27577
rect 522 27521 590 27577
rect 646 27521 714 27577
rect 770 27521 838 27577
rect 894 27521 1000 27577
rect 0 27453 1000 27521
rect 0 27397 94 27453
rect 150 27397 218 27453
rect 274 27397 342 27453
rect 398 27397 466 27453
rect 522 27397 590 27453
rect 646 27397 714 27453
rect 770 27397 838 27453
rect 894 27397 1000 27453
rect 0 27329 1000 27397
rect 0 27273 94 27329
rect 150 27273 218 27329
rect 274 27273 342 27329
rect 398 27273 466 27329
rect 522 27273 590 27329
rect 646 27273 714 27329
rect 770 27273 838 27329
rect 894 27273 1000 27329
rect 0 27205 1000 27273
rect 0 27149 94 27205
rect 150 27149 218 27205
rect 274 27149 342 27205
rect 398 27149 466 27205
rect 522 27149 590 27205
rect 646 27149 714 27205
rect 770 27149 838 27205
rect 894 27149 1000 27205
rect 0 27081 1000 27149
rect 0 27025 94 27081
rect 150 27025 218 27081
rect 274 27025 342 27081
rect 398 27025 466 27081
rect 522 27025 590 27081
rect 646 27025 714 27081
rect 770 27025 838 27081
rect 894 27025 1000 27081
rect 0 26957 1000 27025
rect 0 26901 94 26957
rect 150 26901 218 26957
rect 274 26901 342 26957
rect 398 26901 466 26957
rect 522 26901 590 26957
rect 646 26901 714 26957
rect 770 26901 838 26957
rect 894 26901 1000 26957
rect 0 26800 1000 26901
rect 0 26496 1000 26600
rect 0 26440 95 26496
rect 151 26440 219 26496
rect 275 26440 343 26496
rect 399 26440 467 26496
rect 523 26440 591 26496
rect 647 26440 715 26496
rect 771 26440 839 26496
rect 895 26440 1000 26496
rect 0 26372 1000 26440
rect 0 26316 95 26372
rect 151 26316 219 26372
rect 275 26316 343 26372
rect 399 26316 467 26372
rect 523 26316 591 26372
rect 647 26316 715 26372
rect 771 26316 839 26372
rect 895 26316 1000 26372
rect 0 26248 1000 26316
rect 0 26192 95 26248
rect 151 26192 219 26248
rect 275 26192 343 26248
rect 399 26192 467 26248
rect 523 26192 591 26248
rect 647 26192 715 26248
rect 771 26192 839 26248
rect 895 26192 1000 26248
rect 0 26124 1000 26192
rect 0 26068 95 26124
rect 151 26068 219 26124
rect 275 26068 343 26124
rect 399 26068 467 26124
rect 523 26068 591 26124
rect 647 26068 715 26124
rect 771 26068 839 26124
rect 895 26068 1000 26124
rect 0 26000 1000 26068
rect 0 25944 95 26000
rect 151 25944 219 26000
rect 275 25944 343 26000
rect 399 25944 467 26000
rect 523 25944 591 26000
rect 647 25944 715 26000
rect 771 25944 839 26000
rect 895 25944 1000 26000
rect 0 25876 1000 25944
rect 0 25820 95 25876
rect 151 25820 219 25876
rect 275 25820 343 25876
rect 399 25820 467 25876
rect 523 25820 591 25876
rect 647 25820 715 25876
rect 771 25820 839 25876
rect 895 25820 1000 25876
rect 0 25752 1000 25820
rect 0 25696 95 25752
rect 151 25696 219 25752
rect 275 25696 343 25752
rect 399 25696 467 25752
rect 523 25696 591 25752
rect 647 25696 715 25752
rect 771 25696 839 25752
rect 895 25696 1000 25752
rect 0 25628 1000 25696
rect 0 25572 95 25628
rect 151 25572 219 25628
rect 275 25572 343 25628
rect 399 25572 467 25628
rect 523 25572 591 25628
rect 647 25572 715 25628
rect 771 25572 839 25628
rect 895 25572 1000 25628
rect 0 25504 1000 25572
rect 0 25448 95 25504
rect 151 25448 219 25504
rect 275 25448 343 25504
rect 399 25448 467 25504
rect 523 25448 591 25504
rect 647 25448 715 25504
rect 771 25448 839 25504
rect 895 25448 1000 25504
rect 0 25380 1000 25448
rect 0 25324 95 25380
rect 151 25324 219 25380
rect 275 25324 343 25380
rect 399 25324 467 25380
rect 523 25324 591 25380
rect 647 25324 715 25380
rect 771 25324 839 25380
rect 895 25324 1000 25380
rect 0 25200 1000 25324
rect 0 24884 1000 25000
rect 0 24828 95 24884
rect 151 24828 219 24884
rect 275 24828 343 24884
rect 399 24828 467 24884
rect 523 24828 591 24884
rect 647 24828 715 24884
rect 771 24828 839 24884
rect 895 24828 1000 24884
rect 0 24760 1000 24828
rect 0 24704 95 24760
rect 151 24704 219 24760
rect 275 24704 343 24760
rect 399 24704 467 24760
rect 523 24704 591 24760
rect 647 24704 715 24760
rect 771 24704 839 24760
rect 895 24704 1000 24760
rect 0 24636 1000 24704
rect 0 24580 95 24636
rect 151 24580 219 24636
rect 275 24580 343 24636
rect 399 24580 467 24636
rect 523 24580 591 24636
rect 647 24580 715 24636
rect 771 24580 839 24636
rect 895 24580 1000 24636
rect 0 24512 1000 24580
rect 0 24456 95 24512
rect 151 24456 219 24512
rect 275 24456 343 24512
rect 399 24456 467 24512
rect 523 24456 591 24512
rect 647 24456 715 24512
rect 771 24456 839 24512
rect 895 24456 1000 24512
rect 0 24388 1000 24456
rect 0 24332 95 24388
rect 151 24332 219 24388
rect 275 24332 343 24388
rect 399 24332 467 24388
rect 523 24332 591 24388
rect 647 24332 715 24388
rect 771 24332 839 24388
rect 895 24332 1000 24388
rect 0 24264 1000 24332
rect 0 24208 95 24264
rect 151 24208 219 24264
rect 275 24208 343 24264
rect 399 24208 467 24264
rect 523 24208 591 24264
rect 647 24208 715 24264
rect 771 24208 839 24264
rect 895 24208 1000 24264
rect 0 24140 1000 24208
rect 0 24084 95 24140
rect 151 24084 219 24140
rect 275 24084 343 24140
rect 399 24084 467 24140
rect 523 24084 591 24140
rect 647 24084 715 24140
rect 771 24084 839 24140
rect 895 24084 1000 24140
rect 0 24016 1000 24084
rect 0 23960 95 24016
rect 151 23960 219 24016
rect 275 23960 343 24016
rect 399 23960 467 24016
rect 523 23960 591 24016
rect 647 23960 715 24016
rect 771 23960 839 24016
rect 895 23960 1000 24016
rect 0 23892 1000 23960
rect 0 23836 95 23892
rect 151 23836 219 23892
rect 275 23836 343 23892
rect 399 23836 467 23892
rect 523 23836 591 23892
rect 647 23836 715 23892
rect 771 23836 839 23892
rect 895 23836 1000 23892
rect 0 23768 1000 23836
rect 0 23712 95 23768
rect 151 23712 219 23768
rect 275 23712 343 23768
rect 399 23712 467 23768
rect 523 23712 591 23768
rect 647 23712 715 23768
rect 771 23712 839 23768
rect 895 23712 1000 23768
rect 0 23600 1000 23712
rect 0 23297 1000 23400
rect 0 23241 94 23297
rect 150 23241 218 23297
rect 274 23241 342 23297
rect 398 23241 466 23297
rect 522 23241 590 23297
rect 646 23241 714 23297
rect 770 23241 838 23297
rect 894 23241 1000 23297
rect 0 23173 1000 23241
rect 0 23117 94 23173
rect 150 23117 218 23173
rect 274 23117 342 23173
rect 398 23117 466 23173
rect 522 23117 590 23173
rect 646 23117 714 23173
rect 770 23117 838 23173
rect 894 23117 1000 23173
rect 0 23049 1000 23117
rect 0 22993 94 23049
rect 150 22993 218 23049
rect 274 22993 342 23049
rect 398 22993 466 23049
rect 522 22993 590 23049
rect 646 22993 714 23049
rect 770 22993 838 23049
rect 894 22993 1000 23049
rect 0 22925 1000 22993
rect 0 22869 94 22925
rect 150 22869 218 22925
rect 274 22869 342 22925
rect 398 22869 466 22925
rect 522 22869 590 22925
rect 646 22869 714 22925
rect 770 22869 838 22925
rect 894 22869 1000 22925
rect 0 22801 1000 22869
rect 0 22745 94 22801
rect 150 22745 218 22801
rect 274 22745 342 22801
rect 398 22745 466 22801
rect 522 22745 590 22801
rect 646 22745 714 22801
rect 770 22745 838 22801
rect 894 22745 1000 22801
rect 0 22677 1000 22745
rect 0 22621 94 22677
rect 150 22621 218 22677
rect 274 22621 342 22677
rect 398 22621 466 22677
rect 522 22621 590 22677
rect 646 22621 714 22677
rect 770 22621 838 22677
rect 894 22621 1000 22677
rect 0 22553 1000 22621
rect 0 22497 94 22553
rect 150 22497 218 22553
rect 274 22497 342 22553
rect 398 22497 466 22553
rect 522 22497 590 22553
rect 646 22497 714 22553
rect 770 22497 838 22553
rect 894 22497 1000 22553
rect 0 22429 1000 22497
rect 0 22373 94 22429
rect 150 22373 218 22429
rect 274 22373 342 22429
rect 398 22373 466 22429
rect 522 22373 590 22429
rect 646 22373 714 22429
rect 770 22373 838 22429
rect 894 22373 1000 22429
rect 0 22305 1000 22373
rect 0 22249 94 22305
rect 150 22249 218 22305
rect 274 22249 342 22305
rect 398 22249 466 22305
rect 522 22249 590 22305
rect 646 22249 714 22305
rect 770 22249 838 22305
rect 894 22249 1000 22305
rect 0 22181 1000 22249
rect 0 22125 94 22181
rect 150 22125 218 22181
rect 274 22125 342 22181
rect 398 22125 466 22181
rect 522 22125 590 22181
rect 646 22125 714 22181
rect 770 22125 838 22181
rect 894 22125 1000 22181
rect 0 22057 1000 22125
rect 0 22001 94 22057
rect 150 22001 218 22057
rect 274 22001 342 22057
rect 398 22001 466 22057
rect 522 22001 590 22057
rect 646 22001 714 22057
rect 770 22001 838 22057
rect 894 22001 1000 22057
rect 0 21933 1000 22001
rect 0 21877 94 21933
rect 150 21877 218 21933
rect 274 21877 342 21933
rect 398 21877 466 21933
rect 522 21877 590 21933
rect 646 21877 714 21933
rect 770 21877 838 21933
rect 894 21877 1000 21933
rect 0 21809 1000 21877
rect 0 21753 94 21809
rect 150 21753 218 21809
rect 274 21753 342 21809
rect 398 21753 466 21809
rect 522 21753 590 21809
rect 646 21753 714 21809
rect 770 21753 838 21809
rect 894 21753 1000 21809
rect 0 21685 1000 21753
rect 0 21629 94 21685
rect 150 21629 218 21685
rect 274 21629 342 21685
rect 398 21629 466 21685
rect 522 21629 590 21685
rect 646 21629 714 21685
rect 770 21629 838 21685
rect 894 21629 1000 21685
rect 0 21561 1000 21629
rect 0 21505 94 21561
rect 150 21505 218 21561
rect 274 21505 342 21561
rect 398 21505 466 21561
rect 522 21505 590 21561
rect 646 21505 714 21561
rect 770 21505 838 21561
rect 894 21505 1000 21561
rect 0 21437 1000 21505
rect 0 21381 94 21437
rect 150 21381 218 21437
rect 274 21381 342 21437
rect 398 21381 466 21437
rect 522 21381 590 21437
rect 646 21381 714 21437
rect 770 21381 838 21437
rect 894 21381 1000 21437
rect 0 21313 1000 21381
rect 0 21257 94 21313
rect 150 21257 218 21313
rect 274 21257 342 21313
rect 398 21257 466 21313
rect 522 21257 590 21313
rect 646 21257 714 21313
rect 770 21257 838 21313
rect 894 21257 1000 21313
rect 0 21189 1000 21257
rect 0 21133 94 21189
rect 150 21133 218 21189
rect 274 21133 342 21189
rect 398 21133 466 21189
rect 522 21133 590 21189
rect 646 21133 714 21189
rect 770 21133 838 21189
rect 894 21133 1000 21189
rect 0 21065 1000 21133
rect 0 21009 94 21065
rect 150 21009 218 21065
rect 274 21009 342 21065
rect 398 21009 466 21065
rect 522 21009 590 21065
rect 646 21009 714 21065
rect 770 21009 838 21065
rect 894 21009 1000 21065
rect 0 20941 1000 21009
rect 0 20885 94 20941
rect 150 20885 218 20941
rect 274 20885 342 20941
rect 398 20885 466 20941
rect 522 20885 590 20941
rect 646 20885 714 20941
rect 770 20885 838 20941
rect 894 20885 1000 20941
rect 0 20817 1000 20885
rect 0 20761 94 20817
rect 150 20761 218 20817
rect 274 20761 342 20817
rect 398 20761 466 20817
rect 522 20761 590 20817
rect 646 20761 714 20817
rect 770 20761 838 20817
rect 894 20761 1000 20817
rect 0 20693 1000 20761
rect 0 20637 94 20693
rect 150 20637 218 20693
rect 274 20637 342 20693
rect 398 20637 466 20693
rect 522 20637 590 20693
rect 646 20637 714 20693
rect 770 20637 838 20693
rect 894 20637 1000 20693
rect 0 20569 1000 20637
rect 0 20513 94 20569
rect 150 20513 218 20569
rect 274 20513 342 20569
rect 398 20513 466 20569
rect 522 20513 590 20569
rect 646 20513 714 20569
rect 770 20513 838 20569
rect 894 20513 1000 20569
rect 0 20400 1000 20513
rect 0 20086 1000 20200
rect 0 20030 94 20086
rect 150 20030 218 20086
rect 274 20030 342 20086
rect 398 20030 466 20086
rect 522 20030 590 20086
rect 646 20030 714 20086
rect 770 20030 838 20086
rect 894 20030 1000 20086
rect 0 19962 1000 20030
rect 0 19906 94 19962
rect 150 19906 218 19962
rect 274 19906 342 19962
rect 398 19906 466 19962
rect 522 19906 590 19962
rect 646 19906 714 19962
rect 770 19906 838 19962
rect 894 19906 1000 19962
rect 0 19838 1000 19906
rect 0 19782 94 19838
rect 150 19782 218 19838
rect 274 19782 342 19838
rect 398 19782 466 19838
rect 522 19782 590 19838
rect 646 19782 714 19838
rect 770 19782 838 19838
rect 894 19782 1000 19838
rect 0 19714 1000 19782
rect 0 19658 94 19714
rect 150 19658 218 19714
rect 274 19658 342 19714
rect 398 19658 466 19714
rect 522 19658 590 19714
rect 646 19658 714 19714
rect 770 19658 838 19714
rect 894 19658 1000 19714
rect 0 19590 1000 19658
rect 0 19534 94 19590
rect 150 19534 218 19590
rect 274 19534 342 19590
rect 398 19534 466 19590
rect 522 19534 590 19590
rect 646 19534 714 19590
rect 770 19534 838 19590
rect 894 19534 1000 19590
rect 0 19466 1000 19534
rect 0 19410 94 19466
rect 150 19410 218 19466
rect 274 19410 342 19466
rect 398 19410 466 19466
rect 522 19410 590 19466
rect 646 19410 714 19466
rect 770 19410 838 19466
rect 894 19410 1000 19466
rect 0 19342 1000 19410
rect 0 19286 94 19342
rect 150 19286 218 19342
rect 274 19286 342 19342
rect 398 19286 466 19342
rect 522 19286 590 19342
rect 646 19286 714 19342
rect 770 19286 838 19342
rect 894 19286 1000 19342
rect 0 19218 1000 19286
rect 0 19162 94 19218
rect 150 19162 218 19218
rect 274 19162 342 19218
rect 398 19162 466 19218
rect 522 19162 590 19218
rect 646 19162 714 19218
rect 770 19162 838 19218
rect 894 19162 1000 19218
rect 0 19094 1000 19162
rect 0 19038 94 19094
rect 150 19038 218 19094
rect 274 19038 342 19094
rect 398 19038 466 19094
rect 522 19038 590 19094
rect 646 19038 714 19094
rect 770 19038 838 19094
rect 894 19038 1000 19094
rect 0 18970 1000 19038
rect 0 18914 94 18970
rect 150 18914 218 18970
rect 274 18914 342 18970
rect 398 18914 466 18970
rect 522 18914 590 18970
rect 646 18914 714 18970
rect 770 18914 838 18970
rect 894 18914 1000 18970
rect 0 18846 1000 18914
rect 0 18790 94 18846
rect 150 18790 218 18846
rect 274 18790 342 18846
rect 398 18790 466 18846
rect 522 18790 590 18846
rect 646 18790 714 18846
rect 770 18790 838 18846
rect 894 18790 1000 18846
rect 0 18722 1000 18790
rect 0 18666 94 18722
rect 150 18666 218 18722
rect 274 18666 342 18722
rect 398 18666 466 18722
rect 522 18666 590 18722
rect 646 18666 714 18722
rect 770 18666 838 18722
rect 894 18666 1000 18722
rect 0 18598 1000 18666
rect 0 18542 94 18598
rect 150 18542 218 18598
rect 274 18542 342 18598
rect 398 18542 466 18598
rect 522 18542 590 18598
rect 646 18542 714 18598
rect 770 18542 838 18598
rect 894 18542 1000 18598
rect 0 18474 1000 18542
rect 0 18418 94 18474
rect 150 18418 218 18474
rect 274 18418 342 18474
rect 398 18418 466 18474
rect 522 18418 590 18474
rect 646 18418 714 18474
rect 770 18418 838 18474
rect 894 18418 1000 18474
rect 0 18350 1000 18418
rect 0 18294 94 18350
rect 150 18294 218 18350
rect 274 18294 342 18350
rect 398 18294 466 18350
rect 522 18294 590 18350
rect 646 18294 714 18350
rect 770 18294 838 18350
rect 894 18294 1000 18350
rect 0 18226 1000 18294
rect 0 18170 94 18226
rect 150 18170 218 18226
rect 274 18170 342 18226
rect 398 18170 466 18226
rect 522 18170 590 18226
rect 646 18170 714 18226
rect 770 18170 838 18226
rect 894 18170 1000 18226
rect 0 18102 1000 18170
rect 0 18046 94 18102
rect 150 18046 218 18102
rect 274 18046 342 18102
rect 398 18046 466 18102
rect 522 18046 590 18102
rect 646 18046 714 18102
rect 770 18046 838 18102
rect 894 18046 1000 18102
rect 0 17978 1000 18046
rect 0 17922 94 17978
rect 150 17922 218 17978
rect 274 17922 342 17978
rect 398 17922 466 17978
rect 522 17922 590 17978
rect 646 17922 714 17978
rect 770 17922 838 17978
rect 894 17922 1000 17978
rect 0 17854 1000 17922
rect 0 17798 94 17854
rect 150 17798 218 17854
rect 274 17798 342 17854
rect 398 17798 466 17854
rect 522 17798 590 17854
rect 646 17798 714 17854
rect 770 17798 838 17854
rect 894 17798 1000 17854
rect 0 17730 1000 17798
rect 0 17674 94 17730
rect 150 17674 218 17730
rect 274 17674 342 17730
rect 398 17674 466 17730
rect 522 17674 590 17730
rect 646 17674 714 17730
rect 770 17674 838 17730
rect 894 17674 1000 17730
rect 0 17606 1000 17674
rect 0 17550 94 17606
rect 150 17550 218 17606
rect 274 17550 342 17606
rect 398 17550 466 17606
rect 522 17550 590 17606
rect 646 17550 714 17606
rect 770 17550 838 17606
rect 894 17550 1000 17606
rect 0 17482 1000 17550
rect 0 17426 94 17482
rect 150 17426 218 17482
rect 274 17426 342 17482
rect 398 17426 466 17482
rect 522 17426 590 17482
rect 646 17426 714 17482
rect 770 17426 838 17482
rect 894 17426 1000 17482
rect 0 17358 1000 17426
rect 0 17302 94 17358
rect 150 17302 218 17358
rect 274 17302 342 17358
rect 398 17302 466 17358
rect 522 17302 590 17358
rect 646 17302 714 17358
rect 770 17302 838 17358
rect 894 17302 1000 17358
rect 0 17200 1000 17302
rect 0 16913 1000 17000
rect 0 16857 94 16913
rect 150 16857 218 16913
rect 274 16857 342 16913
rect 398 16857 466 16913
rect 522 16857 590 16913
rect 646 16857 714 16913
rect 770 16857 838 16913
rect 894 16857 1000 16913
rect 0 16789 1000 16857
rect 0 16733 94 16789
rect 150 16733 218 16789
rect 274 16733 342 16789
rect 398 16733 466 16789
rect 522 16733 590 16789
rect 646 16733 714 16789
rect 770 16733 838 16789
rect 894 16733 1000 16789
rect 0 16665 1000 16733
rect 0 16609 94 16665
rect 150 16609 218 16665
rect 274 16609 342 16665
rect 398 16609 466 16665
rect 522 16609 590 16665
rect 646 16609 714 16665
rect 770 16609 838 16665
rect 894 16609 1000 16665
rect 0 16541 1000 16609
rect 0 16485 94 16541
rect 150 16485 218 16541
rect 274 16485 342 16541
rect 398 16485 466 16541
rect 522 16485 590 16541
rect 646 16485 714 16541
rect 770 16485 838 16541
rect 894 16485 1000 16541
rect 0 16417 1000 16485
rect 0 16361 94 16417
rect 150 16361 218 16417
rect 274 16361 342 16417
rect 398 16361 466 16417
rect 522 16361 590 16417
rect 646 16361 714 16417
rect 770 16361 838 16417
rect 894 16361 1000 16417
rect 0 16293 1000 16361
rect 0 16237 94 16293
rect 150 16237 218 16293
rect 274 16237 342 16293
rect 398 16237 466 16293
rect 522 16237 590 16293
rect 646 16237 714 16293
rect 770 16237 838 16293
rect 894 16237 1000 16293
rect 0 16169 1000 16237
rect 0 16113 94 16169
rect 150 16113 218 16169
rect 274 16113 342 16169
rect 398 16113 466 16169
rect 522 16113 590 16169
rect 646 16113 714 16169
rect 770 16113 838 16169
rect 894 16113 1000 16169
rect 0 16045 1000 16113
rect 0 15989 94 16045
rect 150 15989 218 16045
rect 274 15989 342 16045
rect 398 15989 466 16045
rect 522 15989 590 16045
rect 646 15989 714 16045
rect 770 15989 838 16045
rect 894 15989 1000 16045
rect 0 15921 1000 15989
rect 0 15865 94 15921
rect 150 15865 218 15921
rect 274 15865 342 15921
rect 398 15865 466 15921
rect 522 15865 590 15921
rect 646 15865 714 15921
rect 770 15865 838 15921
rect 894 15865 1000 15921
rect 0 15797 1000 15865
rect 0 15741 94 15797
rect 150 15741 218 15797
rect 274 15741 342 15797
rect 398 15741 466 15797
rect 522 15741 590 15797
rect 646 15741 714 15797
rect 770 15741 838 15797
rect 894 15741 1000 15797
rect 0 15673 1000 15741
rect 0 15617 94 15673
rect 150 15617 218 15673
rect 274 15617 342 15673
rect 398 15617 466 15673
rect 522 15617 590 15673
rect 646 15617 714 15673
rect 770 15617 838 15673
rect 894 15617 1000 15673
rect 0 15549 1000 15617
rect 0 15493 94 15549
rect 150 15493 218 15549
rect 274 15493 342 15549
rect 398 15493 466 15549
rect 522 15493 590 15549
rect 646 15493 714 15549
rect 770 15493 838 15549
rect 894 15493 1000 15549
rect 0 15425 1000 15493
rect 0 15369 94 15425
rect 150 15369 218 15425
rect 274 15369 342 15425
rect 398 15369 466 15425
rect 522 15369 590 15425
rect 646 15369 714 15425
rect 770 15369 838 15425
rect 894 15369 1000 15425
rect 0 15301 1000 15369
rect 0 15245 94 15301
rect 150 15245 218 15301
rect 274 15245 342 15301
rect 398 15245 466 15301
rect 522 15245 590 15301
rect 646 15245 714 15301
rect 770 15245 838 15301
rect 894 15245 1000 15301
rect 0 15177 1000 15245
rect 0 15121 94 15177
rect 150 15121 218 15177
rect 274 15121 342 15177
rect 398 15121 466 15177
rect 522 15121 590 15177
rect 646 15121 714 15177
rect 770 15121 838 15177
rect 894 15121 1000 15177
rect 0 15053 1000 15121
rect 0 14997 94 15053
rect 150 14997 218 15053
rect 274 14997 342 15053
rect 398 14997 466 15053
rect 522 14997 590 15053
rect 646 14997 714 15053
rect 770 14997 838 15053
rect 894 14997 1000 15053
rect 0 14929 1000 14997
rect 0 14873 94 14929
rect 150 14873 218 14929
rect 274 14873 342 14929
rect 398 14873 466 14929
rect 522 14873 590 14929
rect 646 14873 714 14929
rect 770 14873 838 14929
rect 894 14873 1000 14929
rect 0 14805 1000 14873
rect 0 14749 94 14805
rect 150 14749 218 14805
rect 274 14749 342 14805
rect 398 14749 466 14805
rect 522 14749 590 14805
rect 646 14749 714 14805
rect 770 14749 838 14805
rect 894 14749 1000 14805
rect 0 14681 1000 14749
rect 0 14625 94 14681
rect 150 14625 218 14681
rect 274 14625 342 14681
rect 398 14625 466 14681
rect 522 14625 590 14681
rect 646 14625 714 14681
rect 770 14625 838 14681
rect 894 14625 1000 14681
rect 0 14557 1000 14625
rect 0 14501 94 14557
rect 150 14501 218 14557
rect 274 14501 342 14557
rect 398 14501 466 14557
rect 522 14501 590 14557
rect 646 14501 714 14557
rect 770 14501 838 14557
rect 894 14501 1000 14557
rect 0 14433 1000 14501
rect 0 14377 94 14433
rect 150 14377 218 14433
rect 274 14377 342 14433
rect 398 14377 466 14433
rect 522 14377 590 14433
rect 646 14377 714 14433
rect 770 14377 838 14433
rect 894 14377 1000 14433
rect 0 14309 1000 14377
rect 0 14253 94 14309
rect 150 14253 218 14309
rect 274 14253 342 14309
rect 398 14253 466 14309
rect 522 14253 590 14309
rect 646 14253 714 14309
rect 770 14253 838 14309
rect 894 14253 1000 14309
rect 0 14185 1000 14253
rect 0 14129 94 14185
rect 150 14129 218 14185
rect 274 14129 342 14185
rect 398 14129 466 14185
rect 522 14129 590 14185
rect 646 14129 714 14185
rect 770 14129 838 14185
rect 894 14129 1000 14185
rect 0 14000 1000 14129
use GF_NI_FILL5_0  GF_NI_FILL5_0_0
timestamp 1666464484
transform 1 0 0 0 1 0
box -32 13097 1032 69968
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_0
timestamp 1666464484
transform 1 0 494 0 1 64300
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_1
timestamp 1666464484
transform 1 0 495 0 1 49894
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_2
timestamp 1666464484
transform 1 0 494 0 1 65891
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_3
timestamp 1666464484
transform 1 0 494 0 1 67498
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_4
timestamp 1666464484
transform 1 0 494 0 1 69043
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_5
timestamp 1666464484
transform 1 0 494 0 1 62694
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_6
timestamp 1666464484
transform 1 0 494 0 1 61108
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_7
timestamp 1666464484
transform 1 0 494 0 1 59516
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_8
timestamp 1666464484
transform 1 0 494 0 1 57899
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_9
timestamp 1666464484
transform 1 0 494 0 1 56306
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_10
timestamp 1666464484
transform 1 0 494 0 1 54702
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_11
timestamp 1666464484
transform 1 0 494 0 1 53096
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_12
timestamp 1666464484
transform 1 0 494 0 1 51493
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_13
timestamp 1666464484
transform 1 0 495 0 1 41898
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_14
timestamp 1666464484
transform 1 0 495 0 1 40310
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_15
timestamp 1666464484
transform 1 0 495 0 1 25910
box 0 0 1 1
use M4_M3_CDNS_40661954729316  M4_M3_CDNS_40661954729316_16
timestamp 1666464484
transform 1 0 495 0 1 24298
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_0
timestamp 1666464484
transform 1 0 494 0 1 44305
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_1
timestamp 1666464484
transform 1 0 494 0 1 37912
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_2
timestamp 1666464484
transform 1 0 494 0 1 34702
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_3
timestamp 1666464484
transform 1 0 494 0 1 31510
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_4
timestamp 1666464484
transform 1 0 494 0 1 28293
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_5
timestamp 1666464484
transform 1 0 494 0 1 21905
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_6
timestamp 1666464484
transform 1 0 494 0 1 18694
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_7
timestamp 1666464484
transform 1 0 494 0 1 15521
box 0 0 1 1
use M4_M3_CDNS_40661954729317  M4_M3_CDNS_40661954729317_8
timestamp 1666464484
transform 1 0 494 0 1 47501
box 0 0 1 1
<< labels >>
rlabel metal4 s 800 14000 1000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 26800 1000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 50800 1000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 800 49200 1000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 800 30000 1000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 17200 1000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 63600 1000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 800 62000 1000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal4 s 800 33200 1000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 36400 1000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 42800 1000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 20400 1000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 23600 1000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 46000 1000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 25200 1000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 39600 1000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 57200 1000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 41200 1000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 60400 1000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 52400 1000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 54000 1000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 55600 1000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 58800 1000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 65200 1000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 800 66800 1000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 800 68400 1000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 26800 1000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 49200 1000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 30000 1000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 33200 1000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 36400 1000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 42800 1000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 23600 1000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 41200 1000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 52400 1000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 54000 1000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 63600 1000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 50800 1000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 62000 1000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 14000 1000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 17200 1000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 20400 1000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 46000 1000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 25200 1000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 39600 1000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 57200 1000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 60400 1000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 65200 1000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 68400 1000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 55600 1000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 58800 1000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 66800 1000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel space 0 400 0 400 4 & Metric 1.00
rlabel space 0 800 0 800 4 & Version 2014q3v1
rlabel space 0 1200 0 1200 4 & Product GF018green_ipio_5p0c_75
rlabel space 0 1600 0 1600 4 & Vendor GLOBALFOUNDRIES
rlabel metal3 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal4 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 68400 200 69678 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 68400 200 69678 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 65200 200 66600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal4 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal4 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 63600 200 65000 1 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 63600 200 65000 1 VSS
port 4 nsew ground bidirectional
rlabel metal4 s 0 49200 200 50600 1 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 1 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string GDS_END 4596436
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4591052
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
