magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 476 2998 1094
rect -86 453 86 476
rect 1813 453 2998 476
<< pwell >>
rect 86 453 1813 476
rect -86 -86 2998 453
<< mvnmos >>
rect 372 284 492 356
rect 124 123 244 195
rect 372 123 492 195
rect 804 261 924 333
rect 1172 261 1292 333
rect 804 117 924 189
rect 1172 117 1292 189
rect 1604 261 1724 333
rect 1604 117 1724 189
rect 1964 69 2084 333
rect 2188 69 2308 333
rect 2412 69 2532 333
rect 2636 69 2756 333
<< mvpmos >>
rect 124 740 224 812
rect 372 740 472 812
rect 372 596 472 668
rect 804 740 904 812
rect 1172 740 1272 812
rect 804 596 904 668
rect 1172 596 1272 668
rect 1604 740 1704 812
rect 1604 596 1704 668
rect 1964 573 2064 939
rect 2188 573 2288 939
rect 2412 573 2512 939
rect 2636 573 2736 939
<< mvndiff >>
rect 284 343 372 356
rect 284 297 297 343
rect 343 297 372 343
rect 284 284 372 297
rect 492 284 612 356
rect 552 195 612 284
rect 36 182 124 195
rect 36 136 49 182
rect 95 136 124 182
rect 36 123 124 136
rect 244 182 372 195
rect 244 136 273 182
rect 319 136 372 182
rect 244 123 372 136
rect 492 123 612 195
rect 684 261 804 333
rect 924 320 1012 333
rect 924 274 953 320
rect 999 274 1012 320
rect 924 261 1012 274
rect 1084 320 1172 333
rect 1084 274 1097 320
rect 1143 274 1172 320
rect 1084 261 1172 274
rect 1292 261 1412 333
rect 684 189 744 261
rect 1352 189 1412 261
rect 684 117 804 189
rect 924 176 1172 189
rect 924 130 953 176
rect 999 130 1172 176
rect 924 117 1172 130
rect 1292 117 1412 189
rect 1484 261 1604 333
rect 1724 320 1812 333
rect 1724 274 1753 320
rect 1799 274 1812 320
rect 1724 261 1812 274
rect 1484 189 1544 261
rect 1884 189 1964 333
rect 1484 117 1604 189
rect 1724 176 1964 189
rect 1724 130 1753 176
rect 1799 130 1964 176
rect 1724 117 1964 130
rect 1884 69 1964 117
rect 2084 320 2188 333
rect 2084 180 2113 320
rect 2159 180 2188 320
rect 2084 69 2188 180
rect 2308 222 2412 333
rect 2308 82 2337 222
rect 2383 82 2412 222
rect 2308 69 2412 82
rect 2532 320 2636 333
rect 2532 180 2561 320
rect 2607 180 2636 320
rect 2532 69 2636 180
rect 2756 222 2844 333
rect 2756 82 2785 222
rect 2831 82 2844 222
rect 2756 69 2844 82
<< mvpdiff >>
rect 1884 812 1964 939
rect 36 799 124 812
rect 36 753 49 799
rect 95 753 124 799
rect 36 740 124 753
rect 224 799 372 812
rect 224 753 253 799
rect 299 753 372 799
rect 224 740 372 753
rect 472 740 592 812
rect 532 668 592 740
rect 284 655 372 668
rect 284 609 297 655
rect 343 609 372 655
rect 284 596 372 609
rect 472 596 592 668
rect 684 740 804 812
rect 904 799 1172 812
rect 904 753 933 799
rect 979 753 1172 799
rect 904 740 1172 753
rect 1272 740 1392 812
rect 684 668 744 740
rect 1332 668 1392 740
rect 684 596 804 668
rect 904 655 992 668
rect 904 609 933 655
rect 979 609 992 655
rect 904 596 992 609
rect 1084 655 1172 668
rect 1084 609 1097 655
rect 1143 609 1172 655
rect 1084 596 1172 609
rect 1272 596 1392 668
rect 1484 740 1604 812
rect 1704 799 1964 812
rect 1704 753 1733 799
rect 1779 753 1964 799
rect 1704 740 1964 753
rect 1484 668 1544 740
rect 1484 596 1604 668
rect 1704 655 1792 668
rect 1704 609 1733 655
rect 1779 609 1792 655
rect 1704 596 1792 609
rect 1884 573 1964 740
rect 2064 726 2188 939
rect 2064 586 2113 726
rect 2159 586 2188 726
rect 2064 573 2188 586
rect 2288 926 2412 939
rect 2288 786 2317 926
rect 2363 786 2412 926
rect 2288 573 2412 786
rect 2512 726 2636 939
rect 2512 586 2541 726
rect 2587 586 2636 726
rect 2512 573 2636 586
rect 2736 926 2824 939
rect 2736 786 2765 926
rect 2811 786 2824 926
rect 2736 573 2824 786
<< mvndiffc >>
rect 297 297 343 343
rect 49 136 95 182
rect 273 136 319 182
rect 953 274 999 320
rect 1097 274 1143 320
rect 953 130 999 176
rect 1753 274 1799 320
rect 1753 130 1799 176
rect 2113 180 2159 320
rect 2337 82 2383 222
rect 2561 180 2607 320
rect 2785 82 2831 222
<< mvpdiffc >>
rect 49 753 95 799
rect 253 753 299 799
rect 297 609 343 655
rect 933 753 979 799
rect 933 609 979 655
rect 1097 609 1143 655
rect 1733 753 1779 799
rect 1733 609 1779 655
rect 2113 586 2159 726
rect 2317 786 2363 926
rect 2541 586 2587 726
rect 2765 786 2811 926
<< polysilicon >>
rect 1964 939 2064 983
rect 2188 939 2288 983
rect 2412 939 2512 983
rect 2636 939 2736 983
rect 124 812 224 856
rect 372 812 472 856
rect 804 812 904 856
rect 1172 812 1272 856
rect 1604 812 1704 856
rect 124 368 224 740
rect 372 668 472 740
rect 804 668 904 740
rect 1172 668 1272 740
rect 1604 668 1704 740
rect 124 228 141 368
rect 187 239 224 368
rect 372 552 472 596
rect 372 412 385 552
rect 431 412 472 552
rect 372 400 472 412
rect 804 506 904 596
rect 372 356 492 400
rect 804 366 817 506
rect 863 377 904 506
rect 1172 506 1272 596
rect 863 366 924 377
rect 804 333 924 366
rect 1172 366 1185 506
rect 1231 377 1272 506
rect 1604 506 1704 596
rect 1231 366 1292 377
rect 1172 333 1292 366
rect 1604 366 1617 506
rect 1663 377 1704 506
rect 1964 465 2064 573
rect 2188 465 2288 573
rect 2412 465 2512 573
rect 2636 465 2736 573
rect 1964 452 2736 465
rect 1964 406 1977 452
rect 2399 406 2736 452
rect 1964 393 2736 406
rect 1663 366 1724 377
rect 1604 333 1724 366
rect 1964 333 2084 393
rect 2188 333 2308 393
rect 2412 333 2532 393
rect 2636 377 2736 393
rect 2636 333 2756 377
rect 187 228 244 239
rect 124 195 244 228
rect 372 195 492 284
rect 804 189 924 261
rect 1172 189 1292 261
rect 124 79 244 123
rect 372 79 492 123
rect 1604 189 1724 261
rect 804 73 924 117
rect 1172 73 1292 117
rect 1604 73 1724 117
rect 1964 25 2084 69
rect 2188 25 2308 69
rect 2412 25 2532 69
rect 2636 25 2756 69
<< polycontact >>
rect 141 228 187 368
rect 385 412 431 552
rect 817 366 863 506
rect 1185 366 1231 506
rect 1617 366 1663 506
rect 1977 406 2399 452
<< metal1 >>
rect 0 926 2912 1098
rect 0 918 2317 926
rect 38 799 95 810
rect 38 753 49 799
rect 38 552 95 753
rect 253 799 299 918
rect 253 742 299 753
rect 933 799 979 918
rect 933 742 979 753
rect 1733 799 1779 918
rect 2363 918 2765 926
rect 2317 775 2363 786
rect 2811 918 2912 926
rect 2765 775 2811 786
rect 1733 742 1779 753
rect 2113 726 2159 737
rect 297 655 863 666
rect 343 609 863 655
rect 297 598 863 609
rect 38 506 385 552
rect 38 182 84 506
rect 374 412 385 506
rect 431 412 442 552
rect 817 506 863 598
rect 130 228 141 368
rect 187 228 198 368
rect 817 343 863 366
rect 286 297 297 343
rect 343 297 863 343
rect 933 655 979 666
rect 933 412 979 609
rect 1097 655 1143 666
rect 1097 598 1143 609
rect 1733 655 1779 666
rect 1097 552 1663 598
rect 1617 506 1663 552
rect 1174 412 1185 506
rect 933 366 1185 412
rect 1231 366 1242 506
rect 933 320 999 366
rect 1617 320 1663 366
rect 933 274 953 320
rect 1086 274 1097 320
rect 1143 274 1663 320
rect 1733 463 1779 609
rect 2541 726 2587 737
rect 2159 586 2541 621
rect 2113 575 2587 586
rect 1733 452 2399 463
rect 1733 406 1977 452
rect 1733 395 2399 406
rect 1733 320 1799 395
rect 2445 331 2491 575
rect 1733 274 1753 320
rect 933 263 999 274
rect 1733 263 1799 274
rect 2113 320 2607 331
rect 273 182 319 193
rect 38 136 49 182
rect 95 136 106 182
rect 273 90 319 136
rect 953 176 999 187
rect 953 90 999 130
rect 1753 176 1799 187
rect 2159 285 2561 320
rect 2113 169 2159 180
rect 2337 222 2383 233
rect 1753 90 1799 130
rect 0 82 2337 90
rect 2494 180 2561 285
rect 2494 169 2607 180
rect 2785 222 2831 233
rect 2383 82 2785 90
rect 2831 82 2912 90
rect 0 -90 2912 82
<< labels >>
flabel metal1 s 130 228 198 368 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 2912 1098 0 FreeSans 200 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 2785 193 2831 233 0 FreeSans 200 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 2541 621 2587 737 0 FreeSans 200 0 0 0 Z
port 2 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 2113 621 2159 737 1 Z
port 2 nsew default output
rlabel metal1 s 2113 575 2587 621 1 Z
port 2 nsew default output
rlabel metal1 s 2445 331 2491 575 1 Z
port 2 nsew default output
rlabel metal1 s 2113 285 2607 331 1 Z
port 2 nsew default output
rlabel metal1 s 2494 169 2607 285 1 Z
port 2 nsew default output
rlabel metal1 s 2113 169 2159 285 1 Z
port 2 nsew default output
rlabel metal1 s 2765 775 2811 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2317 775 2363 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1733 775 1779 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 933 775 979 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 253 775 299 918 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1733 742 1779 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 933 742 979 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 253 742 299 775 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2337 193 2383 233 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2785 187 2831 193 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2337 187 2383 193 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 187 319 193 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2785 90 2831 187 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2337 90 2383 187 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1753 90 1799 187 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 953 90 999 187 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 187 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2912 90 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2912 1008
string GDS_END 726760
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 720034
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
