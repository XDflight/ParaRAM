magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 568 1048
<< polysilicon >>
rect -30 907 88 979
rect 194 907 312 979
rect -30 -74 88 -1
rect 194 -74 312 -1
use pmos_5p04310589983262_64x8m81  pmos_5p04310589983262_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 552 1028
<< properties >>
string GDS_END 50608
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 50166
<< end >>
