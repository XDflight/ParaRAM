magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 5910 1094
<< pwell >>
rect -86 -86 5910 453
<< mvnmos >>
rect 124 199 244 317
rect 348 199 468 317
rect 516 199 636 317
rect 740 199 860 317
rect 908 199 1028 317
rect 1343 175 1463 333
rect 1567 175 1687 333
rect 1951 215 2071 333
rect 2175 215 2295 333
rect 2343 215 2463 333
rect 2543 215 2663 333
rect 2811 215 2931 333
rect 2979 215 3099 333
rect 3203 215 3323 333
rect 3427 215 3547 333
rect 3881 181 4001 299
rect 4049 181 4169 299
rect 4273 181 4393 299
rect 4533 69 4653 333
rect 4901 69 5021 333
rect 5125 69 5245 333
rect 5349 69 5469 333
rect 5573 69 5693 333
<< mvpmos >>
rect 124 652 224 852
rect 328 652 428 852
rect 476 652 576 852
rect 680 652 780 852
rect 828 652 928 852
rect 1215 596 1315 872
rect 1507 596 1607 872
rect 1855 577 1955 777
rect 2059 577 2159 777
rect 2263 577 2363 777
rect 2543 686 2643 886
rect 2891 686 2991 886
rect 3197 577 3297 777
rect 3401 577 3501 777
rect 3605 577 3705 777
rect 3953 667 4053 867
rect 4157 667 4257 867
rect 4405 573 4505 939
rect 4613 573 4713 939
rect 4841 573 4941 939
rect 5045 573 5145 939
rect 5249 573 5349 939
rect 5453 573 5553 939
<< mvndiff >>
rect 36 296 124 317
rect 36 250 49 296
rect 95 250 124 296
rect 36 199 124 250
rect 244 296 348 317
rect 244 250 273 296
rect 319 250 348 296
rect 244 199 348 250
rect 468 199 516 317
rect 636 296 740 317
rect 636 250 665 296
rect 711 250 740 296
rect 636 199 740 250
rect 860 199 908 317
rect 1028 199 1148 317
rect 1088 108 1148 199
rect 1255 301 1343 333
rect 1255 255 1268 301
rect 1314 255 1343 301
rect 1255 175 1343 255
rect 1463 265 1567 333
rect 1463 219 1492 265
rect 1538 219 1567 265
rect 1463 175 1567 219
rect 1687 301 1775 333
rect 1687 255 1716 301
rect 1762 255 1775 301
rect 1687 175 1775 255
rect 1863 296 1951 333
rect 1863 250 1876 296
rect 1922 250 1951 296
rect 1863 215 1951 250
rect 2071 296 2175 333
rect 2071 250 2100 296
rect 2146 250 2175 296
rect 2071 215 2175 250
rect 2295 215 2343 333
rect 2463 215 2543 333
rect 2663 296 2811 333
rect 2663 250 2692 296
rect 2738 250 2811 296
rect 2663 215 2811 250
rect 2931 215 2979 333
rect 3099 296 3203 333
rect 3099 250 3128 296
rect 3174 250 3203 296
rect 3099 215 3203 250
rect 3323 296 3427 333
rect 3323 250 3352 296
rect 3398 250 3427 296
rect 3323 215 3427 250
rect 3547 296 3635 333
rect 4453 299 4533 333
rect 3547 250 3576 296
rect 3622 250 3635 296
rect 3547 215 3635 250
rect 3793 286 3881 299
rect 3793 240 3806 286
rect 3852 240 3881 286
rect 1076 95 1148 108
rect 1076 49 1089 95
rect 1135 49 1148 95
rect 1076 36 1148 49
rect 3793 181 3881 240
rect 4001 181 4049 299
rect 4169 240 4273 299
rect 4169 194 4198 240
rect 4244 194 4273 240
rect 4169 181 4273 194
rect 4393 181 4533 299
rect 4453 69 4533 181
rect 4653 320 4741 333
rect 4653 180 4682 320
rect 4728 180 4741 320
rect 4653 69 4741 180
rect 4813 294 4901 333
rect 4813 154 4826 294
rect 4872 154 4901 294
rect 4813 69 4901 154
rect 5021 320 5125 333
rect 5021 180 5050 320
rect 5096 180 5125 320
rect 5021 69 5125 180
rect 5245 319 5349 333
rect 5245 179 5274 319
rect 5320 179 5349 319
rect 5245 69 5349 179
rect 5469 320 5573 333
rect 5469 180 5498 320
rect 5544 180 5573 320
rect 5469 69 5573 180
rect 5693 319 5781 333
rect 5693 179 5722 319
rect 5768 179 5781 319
rect 5693 69 5781 179
<< mvpdiff >>
rect 988 958 1060 971
rect 988 912 1001 958
rect 1047 912 1060 958
rect 1375 958 1447 971
rect 988 899 1060 912
rect 988 852 1048 899
rect 1375 912 1388 958
rect 1434 912 1447 958
rect 1375 872 1447 912
rect 2411 959 2483 972
rect 2411 913 2424 959
rect 2470 913 2483 959
rect 3051 959 3123 972
rect 36 839 124 852
rect 36 699 49 839
rect 95 699 124 839
rect 36 652 124 699
rect 224 839 328 852
rect 224 699 253 839
rect 299 699 328 839
rect 224 652 328 699
rect 428 652 476 852
rect 576 839 680 852
rect 576 699 605 839
rect 651 699 680 839
rect 576 652 680 699
rect 780 652 828 852
rect 928 652 1048 852
rect 1127 757 1215 872
rect 1127 711 1140 757
rect 1186 711 1215 757
rect 1127 596 1215 711
rect 1315 596 1507 872
rect 1607 763 1695 872
rect 2411 900 2483 913
rect 2423 886 2483 900
rect 3051 913 3064 959
rect 3110 913 3123 959
rect 3051 886 3123 913
rect 2423 777 2543 886
rect 1607 623 1636 763
rect 1682 623 1695 763
rect 1607 596 1695 623
rect 1767 764 1855 777
rect 1767 624 1780 764
rect 1826 624 1855 764
rect 1767 577 1855 624
rect 1955 764 2059 777
rect 1955 624 1984 764
rect 2030 624 2059 764
rect 1955 577 2059 624
rect 2159 745 2263 777
rect 2159 699 2188 745
rect 2234 699 2263 745
rect 2159 577 2263 699
rect 2363 686 2543 777
rect 2643 745 2731 886
rect 2643 699 2672 745
rect 2718 699 2731 745
rect 2643 686 2731 699
rect 2803 745 2891 886
rect 2803 699 2816 745
rect 2862 699 2891 745
rect 2803 686 2891 699
rect 2991 777 3123 886
rect 4317 921 4405 939
rect 4317 875 4330 921
rect 4376 875 4405 921
rect 4317 867 4405 875
rect 3865 854 3953 867
rect 3865 808 3878 854
rect 3924 808 3953 854
rect 2991 686 3197 777
rect 2363 577 2443 686
rect 3117 577 3197 686
rect 3297 745 3401 777
rect 3297 699 3326 745
rect 3372 699 3401 745
rect 3297 577 3401 699
rect 3501 740 3605 777
rect 3501 600 3530 740
rect 3576 600 3605 740
rect 3501 577 3605 600
rect 3705 648 3793 777
rect 3865 667 3953 808
rect 4053 726 4157 867
rect 4053 680 4082 726
rect 4128 680 4157 726
rect 4053 667 4157 680
rect 4257 667 4405 867
rect 3705 602 3734 648
rect 3780 602 3793 648
rect 3705 577 3793 602
rect 4325 573 4405 667
rect 4505 726 4613 939
rect 4505 586 4534 726
rect 4580 586 4613 726
rect 4505 573 4613 586
rect 4713 839 4841 939
rect 4713 699 4742 839
rect 4788 699 4841 839
rect 4713 573 4841 699
rect 4941 839 5045 939
rect 4941 699 4970 839
rect 5016 699 5045 839
rect 4941 573 5045 699
rect 5145 839 5249 939
rect 5145 699 5174 839
rect 5220 699 5249 839
rect 5145 573 5249 699
rect 5349 839 5453 939
rect 5349 699 5378 839
rect 5424 699 5453 839
rect 5349 573 5453 699
rect 5553 839 5641 939
rect 5553 699 5582 839
rect 5628 699 5641 839
rect 5553 573 5641 699
<< mvndiffc >>
rect 49 250 95 296
rect 273 250 319 296
rect 665 250 711 296
rect 1268 255 1314 301
rect 1492 219 1538 265
rect 1716 255 1762 301
rect 1876 250 1922 296
rect 2100 250 2146 296
rect 2692 250 2738 296
rect 3128 250 3174 296
rect 3352 250 3398 296
rect 3576 250 3622 296
rect 3806 240 3852 286
rect 1089 49 1135 95
rect 4198 194 4244 240
rect 4682 180 4728 320
rect 4826 154 4872 294
rect 5050 180 5096 320
rect 5274 179 5320 319
rect 5498 180 5544 320
rect 5722 179 5768 319
<< mvpdiffc >>
rect 1001 912 1047 958
rect 1388 912 1434 958
rect 2424 913 2470 959
rect 49 699 95 839
rect 253 699 299 839
rect 605 699 651 839
rect 1140 711 1186 757
rect 3064 913 3110 959
rect 1636 623 1682 763
rect 1780 624 1826 764
rect 1984 624 2030 764
rect 2188 699 2234 745
rect 2672 699 2718 745
rect 2816 699 2862 745
rect 4330 875 4376 921
rect 3878 808 3924 854
rect 3326 699 3372 745
rect 3530 600 3576 740
rect 4082 680 4128 726
rect 3734 602 3780 648
rect 4534 586 4580 726
rect 4742 699 4788 839
rect 4970 699 5016 839
rect 5174 699 5220 839
rect 5378 699 5424 839
rect 5582 699 5628 839
<< polysilicon >>
rect 124 944 928 984
rect 124 852 224 944
rect 328 852 428 896
rect 476 852 576 896
rect 680 852 780 896
rect 828 852 928 944
rect 1215 872 1315 916
rect 1507 944 1855 984
rect 1507 872 1607 944
rect 1755 909 1855 944
rect 124 500 224 652
rect 328 608 428 652
rect 124 454 137 500
rect 183 454 224 500
rect 124 361 224 454
rect 348 500 428 608
rect 348 454 361 500
rect 407 454 428 500
rect 348 361 428 454
rect 476 500 576 652
rect 476 454 489 500
rect 535 454 576 500
rect 476 441 576 454
rect 680 500 780 652
rect 828 608 928 652
rect 1755 869 2159 909
rect 2059 856 2159 869
rect 1855 777 1955 821
rect 2059 810 2100 856
rect 2146 810 2159 856
rect 2543 886 2643 930
rect 2891 886 2991 930
rect 2059 777 2159 810
rect 2263 777 2363 821
rect 1215 563 1315 596
rect 1215 517 1256 563
rect 1302 517 1315 563
rect 680 454 702 500
rect 748 454 780 500
rect 680 441 780 454
rect 740 361 780 441
rect 908 500 1028 513
rect 908 454 921 500
rect 967 454 1028 500
rect 124 317 244 361
rect 348 317 468 361
rect 516 317 636 361
rect 740 317 860 361
rect 908 317 1028 454
rect 1215 465 1315 517
rect 1507 500 1607 596
rect 3197 944 4053 984
rect 3197 777 3297 944
rect 3401 856 3501 869
rect 3953 867 4053 944
rect 4405 939 4505 983
rect 4613 939 4713 983
rect 4841 939 4941 983
rect 5045 939 5145 983
rect 5249 939 5349 983
rect 5453 939 5553 983
rect 4157 867 4257 911
rect 3401 810 3414 856
rect 3460 810 3501 856
rect 3401 777 3501 810
rect 3605 777 3705 821
rect 1215 393 1443 465
rect 1507 454 1520 500
rect 1566 454 1607 500
rect 1507 441 1607 454
rect 1343 377 1443 393
rect 1567 377 1607 441
rect 1855 500 1955 577
rect 2059 533 2159 577
rect 2263 533 2363 577
rect 1855 454 1868 500
rect 1914 465 1955 500
rect 2323 515 2363 533
rect 2323 502 2463 515
rect 1914 454 2275 465
rect 1855 425 2275 454
rect 2323 456 2384 502
rect 2430 456 2463 502
rect 2323 445 2463 456
rect 2175 412 2275 425
rect 1343 333 1463 377
rect 1567 333 1687 377
rect 1951 333 2071 377
rect 2175 366 2216 412
rect 2262 377 2275 412
rect 2262 366 2295 377
rect 2175 333 2295 366
rect 2343 333 2463 445
rect 2543 377 2643 686
rect 2891 653 2991 686
rect 2891 607 2904 653
rect 2950 607 2991 653
rect 2891 594 2991 607
rect 2891 377 2931 594
rect 3953 607 4053 667
rect 3881 594 4053 607
rect 3197 497 3297 577
rect 3401 533 3501 577
rect 3605 533 3705 577
rect 2543 333 2663 377
rect 2811 333 2931 377
rect 2979 425 3297 497
rect 2979 333 3099 425
rect 3427 377 3501 533
rect 3665 457 3705 533
rect 3881 548 3942 594
rect 3988 553 4053 594
rect 4157 623 4257 667
rect 3988 548 4001 553
rect 3665 444 3765 457
rect 3665 398 3679 444
rect 3725 398 3765 444
rect 3665 385 3765 398
rect 3203 333 3323 377
rect 3427 333 3547 377
rect 124 107 244 199
rect 348 155 468 199
rect 516 107 636 199
rect 740 155 860 199
rect 908 155 1028 199
rect 3881 299 4001 548
rect 4157 434 4229 623
rect 4405 513 4505 573
rect 4049 422 4229 434
rect 4049 376 4170 422
rect 4216 376 4229 422
rect 4049 363 4229 376
rect 4279 500 4505 513
rect 4279 454 4292 500
rect 4338 473 4505 500
rect 4613 500 4713 573
rect 4338 454 4393 473
rect 4049 299 4169 363
rect 4279 343 4393 454
rect 4613 454 4626 500
rect 4672 454 4713 500
rect 4613 453 4713 454
rect 4553 393 4713 453
rect 4841 513 4941 573
rect 5045 513 5145 573
rect 5249 513 5349 573
rect 5453 513 5553 573
rect 4841 500 5693 513
rect 4841 454 4914 500
rect 4960 454 5693 500
rect 4841 440 5693 454
rect 4553 377 4653 393
rect 4273 299 4393 343
rect 4533 333 4653 377
rect 4901 333 5021 440
rect 5125 333 5245 440
rect 5349 333 5469 440
rect 5573 333 5693 440
rect 1343 131 1463 175
rect 124 35 636 107
rect 1567 107 1687 175
rect 1951 107 2071 215
rect 2175 171 2295 215
rect 2343 171 2463 215
rect 1567 35 2071 107
rect 2543 75 2663 215
rect 2811 171 2931 215
rect 2979 171 3099 215
rect 3203 182 3323 215
rect 3203 136 3216 182
rect 3262 136 3323 182
rect 3427 171 3547 215
rect 3881 137 4001 181
rect 4049 137 4169 181
rect 3203 123 3323 136
rect 4273 75 4393 181
rect 2543 35 4393 75
rect 4533 25 4653 69
rect 4901 25 5021 69
rect 5125 25 5245 69
rect 5349 25 5469 69
rect 5573 25 5693 69
<< polycontact >>
rect 137 454 183 500
rect 361 454 407 500
rect 489 454 535 500
rect 2100 810 2146 856
rect 1256 517 1302 563
rect 702 454 748 500
rect 921 454 967 500
rect 3414 810 3460 856
rect 1520 454 1566 500
rect 1868 454 1914 500
rect 2384 456 2430 502
rect 2216 366 2262 412
rect 2904 607 2950 653
rect 3942 548 3988 594
rect 3679 398 3725 444
rect 4170 376 4216 422
rect 4292 454 4338 500
rect 4626 454 4672 500
rect 4914 454 4960 500
rect 3216 136 3262 182
<< metal1 >>
rect 0 959 5824 1098
rect 0 958 2424 959
rect 0 918 1001 958
rect 49 839 95 850
rect 49 634 95 699
rect 253 839 299 918
rect 990 912 1001 918
rect 1047 918 1388 958
rect 1047 912 1058 918
rect 1377 912 1388 918
rect 1434 918 2424 958
rect 1434 912 1445 918
rect 2470 918 3064 959
rect 2424 902 2470 913
rect 3110 921 5824 959
rect 3110 918 4330 921
rect 3064 902 3110 913
rect 253 688 299 699
rect 605 839 1826 866
rect 651 820 1826 839
rect 1140 757 1566 768
rect 1186 711 1566 757
rect 1140 700 1566 711
rect 605 688 651 699
rect 49 588 967 634
rect 30 500 194 542
rect 30 454 137 500
rect 183 454 194 500
rect 254 500 418 542
rect 254 454 361 500
rect 407 454 418 500
rect 489 500 535 588
rect 489 408 535 454
rect 49 362 535 408
rect 702 500 754 542
rect 748 454 754 500
rect 49 296 95 362
rect 702 354 754 454
rect 921 500 967 588
rect 1150 578 1314 654
rect 1256 563 1314 578
rect 1302 517 1314 563
rect 1256 506 1314 517
rect 1520 500 1566 700
rect 921 443 967 454
rect 1268 454 1520 460
rect 1636 763 1682 774
rect 1636 511 1682 623
rect 1780 764 1826 820
rect 2089 810 2100 856
rect 2146 810 3414 856
rect 3460 810 3471 856
rect 3878 854 3924 918
rect 4319 875 4330 918
rect 4376 918 5824 921
rect 4376 875 4387 918
rect 4742 839 4788 918
rect 3878 797 3924 808
rect 3970 783 4672 829
rect 1780 613 1826 624
rect 1984 764 2030 775
rect 2188 745 2718 756
rect 2234 699 2672 745
rect 2188 688 2718 699
rect 2816 745 3372 756
rect 3970 751 4016 783
rect 2862 710 3326 745
rect 2816 688 2862 699
rect 3128 699 3326 710
rect 3128 688 3372 699
rect 3530 740 4016 751
rect 2904 653 2950 664
rect 2030 642 2110 643
rect 2030 624 2904 642
rect 1984 607 2904 624
rect 1984 597 2950 607
rect 2100 596 2950 597
rect 1636 500 1914 511
rect 1636 465 1868 500
rect 1268 414 1566 454
rect 1716 454 1868 465
rect 1716 443 1914 454
rect 49 239 95 250
rect 273 296 319 307
rect 273 90 319 250
rect 665 296 711 307
rect 665 198 711 250
rect 1268 301 1314 414
rect 1268 244 1314 255
rect 1360 322 1670 368
rect 1360 198 1406 322
rect 665 152 1406 198
rect 1492 265 1538 276
rect 1089 95 1135 106
rect 0 49 1089 90
rect 1492 90 1538 219
rect 1624 198 1670 322
rect 1716 301 1762 443
rect 1716 244 1762 255
rect 1876 296 1922 307
rect 1876 198 1922 250
rect 2100 296 2146 596
rect 3128 513 3174 688
rect 2384 502 3174 513
rect 2430 456 3174 502
rect 2384 445 3174 456
rect 2216 412 2262 423
rect 2262 366 3082 399
rect 2216 353 3082 366
rect 2100 239 2146 250
rect 2692 296 2738 307
rect 1624 152 1922 198
rect 2692 90 2738 250
rect 3036 182 3082 353
rect 3128 296 3174 445
rect 3128 239 3174 250
rect 3352 600 3530 635
rect 3576 705 4016 740
rect 4082 726 4128 737
rect 3352 589 3576 600
rect 3734 648 3780 659
rect 3352 296 3398 589
rect 3734 536 3780 602
rect 3826 594 4002 654
rect 3826 590 3942 594
rect 3931 548 3942 590
rect 3988 548 4002 594
rect 3352 239 3398 250
rect 3576 502 3851 536
rect 4082 502 4128 680
rect 4534 726 4580 737
rect 3576 490 4128 502
rect 3576 296 3622 490
rect 3806 456 4128 490
rect 4286 500 4338 654
rect 3576 239 3622 250
rect 3668 398 3679 444
rect 3725 398 3736 444
rect 3668 182 3736 398
rect 3806 286 3852 456
rect 4286 454 4292 500
rect 4286 443 4338 454
rect 4159 376 4170 422
rect 4216 397 4227 422
rect 4534 397 4580 586
rect 4626 500 4672 783
rect 4742 688 4788 699
rect 4970 839 5016 850
rect 4970 624 5016 699
rect 5174 839 5220 918
rect 5174 688 5220 699
rect 5294 839 5424 850
rect 5294 699 5378 839
rect 5294 688 5424 699
rect 5582 839 5628 918
rect 5582 688 5628 699
rect 5294 624 5346 688
rect 4970 578 5544 624
rect 4626 443 4672 454
rect 4914 500 4960 511
rect 4914 397 4960 454
rect 4216 376 4960 397
rect 4159 351 4960 376
rect 4682 320 4728 351
rect 3806 229 3852 240
rect 4198 240 4244 251
rect 3036 136 3216 182
rect 3262 136 3736 182
rect 4198 90 4244 194
rect 5050 320 5096 578
rect 4682 169 4728 180
rect 4826 294 4872 305
rect 5050 169 5096 180
rect 5274 319 5320 330
rect 4826 90 4872 154
rect 5274 90 5320 179
rect 5498 320 5544 578
rect 5498 169 5544 180
rect 5722 319 5768 330
rect 5722 90 5768 179
rect 1135 49 5824 90
rect 0 -90 5824 49
<< labels >>
flabel metal1 s 1150 578 1314 654 0 FreeSans 200 0 0 0 CLK
port 6 nsew clock input
flabel metal1 s 702 354 754 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 5294 688 5424 850 0 FreeSans 200 0 0 0 Q
port 7 nsew default output
flabel metal1 s 4286 443 4338 654 0 FreeSans 200 0 0 0 RN
port 2 nsew default input
flabel metal1 s 30 454 194 542 0 FreeSans 200 0 0 0 SE
port 3 nsew default input
flabel metal1 s 3826 590 4002 654 0 FreeSans 200 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 254 454 418 542 0 FreeSans 200 0 0 0 SI
port 5 nsew default input
flabel metal1 s 0 918 5824 1098 0 FreeSans 200 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 5722 307 5768 330 0 FreeSans 200 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3931 548 4002 590 1 SETN
port 4 nsew default input
rlabel metal1 s 1256 506 1314 578 1 CLK
port 6 nsew clock input
rlabel metal1 s 4970 688 5016 850 1 Q
port 7 nsew default output
rlabel metal1 s 5294 624 5346 688 1 Q
port 7 nsew default output
rlabel metal1 s 4970 624 5016 688 1 Q
port 7 nsew default output
rlabel metal1 s 4970 578 5544 624 1 Q
port 7 nsew default output
rlabel metal1 s 5498 169 5544 578 1 Q
port 7 nsew default output
rlabel metal1 s 5050 169 5096 578 1 Q
port 7 nsew default output
rlabel metal1 s 5582 912 5628 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5174 912 5220 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4742 912 4788 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4319 912 4387 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3878 912 3924 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3064 912 3110 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2424 912 2470 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1377 912 1445 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 990 912 1058 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 253 912 299 918 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5582 902 5628 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5174 902 5220 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4742 902 4788 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4319 902 4387 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3878 902 3924 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3064 902 3110 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2424 902 2470 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 253 902 299 912 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5582 875 5628 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5174 875 5220 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4742 875 4788 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4319 875 4387 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3878 875 3924 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 253 875 299 902 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5582 797 5628 875 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5174 797 5220 875 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4742 797 4788 875 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3878 797 3924 875 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 253 797 299 875 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5582 688 5628 797 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5174 688 5220 797 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4742 688 4788 797 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 253 688 299 797 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5274 307 5320 330 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5722 305 5768 307 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5274 305 5320 307 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2692 305 2738 307 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 305 319 307 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5722 276 5768 305 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5274 276 5320 305 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4826 276 4872 305 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2692 276 2738 305 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 276 319 305 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5722 251 5768 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5274 251 5320 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4826 251 4872 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2692 251 2738 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1492 251 1538 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 251 319 276 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5722 106 5768 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5274 106 5320 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4826 106 4872 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4198 106 4244 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2692 106 2738 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1492 106 1538 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 106 319 251 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5722 90 5768 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5274 90 5320 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4826 90 4872 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4198 90 4244 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2692 90 2738 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1492 90 1538 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1089 90 1135 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 106 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 5824 90 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5824 1008
string GDS_END 397032
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 384120
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
