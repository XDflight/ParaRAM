magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -19 540 19 546
rect -19 514 -13 540
rect 13 514 19 540
rect -19 478 19 514
rect -19 452 -13 478
rect 13 452 19 478
rect -19 416 19 452
rect -19 390 -13 416
rect 13 390 19 416
rect -19 354 19 390
rect -19 328 -13 354
rect 13 328 19 354
rect -19 292 19 328
rect -19 266 -13 292
rect 13 266 19 292
rect -19 230 19 266
rect -19 204 -13 230
rect 13 204 19 230
rect -19 168 19 204
rect -19 142 -13 168
rect 13 142 19 168
rect -19 106 19 142
rect -19 80 -13 106
rect 13 80 19 106
rect -19 44 19 80
rect -19 18 -13 44
rect 13 18 19 44
rect -19 -18 19 18
rect -19 -44 -13 -18
rect 13 -44 19 -18
rect -19 -80 19 -44
rect -19 -106 -13 -80
rect 13 -106 19 -80
rect -19 -142 19 -106
rect -19 -168 -13 -142
rect 13 -168 19 -142
rect -19 -204 19 -168
rect -19 -230 -13 -204
rect 13 -230 19 -204
rect -19 -266 19 -230
rect -19 -292 -13 -266
rect 13 -292 19 -266
rect -19 -328 19 -292
rect -19 -354 -13 -328
rect 13 -354 19 -328
rect -19 -390 19 -354
rect -19 -416 -13 -390
rect 13 -416 19 -390
rect -19 -452 19 -416
rect -19 -478 -13 -452
rect 13 -478 19 -452
rect -19 -514 19 -478
rect -19 -540 -13 -514
rect 13 -540 19 -514
rect -19 -546 19 -540
<< via1 >>
rect -13 514 13 540
rect -13 452 13 478
rect -13 390 13 416
rect -13 328 13 354
rect -13 266 13 292
rect -13 204 13 230
rect -13 142 13 168
rect -13 80 13 106
rect -13 18 13 44
rect -13 -44 13 -18
rect -13 -106 13 -80
rect -13 -168 13 -142
rect -13 -230 13 -204
rect -13 -292 13 -266
rect -13 -354 13 -328
rect -13 -416 13 -390
rect -13 -478 13 -452
rect -13 -540 13 -514
<< metal2 >>
rect -19 540 19 546
rect -19 514 -13 540
rect 13 514 19 540
rect -19 478 19 514
rect -19 452 -13 478
rect 13 452 19 478
rect -19 416 19 452
rect -19 390 -13 416
rect 13 390 19 416
rect -19 354 19 390
rect -19 328 -13 354
rect 13 328 19 354
rect -19 292 19 328
rect -19 266 -13 292
rect 13 266 19 292
rect -19 230 19 266
rect -19 204 -13 230
rect 13 204 19 230
rect -19 168 19 204
rect -19 142 -13 168
rect 13 142 19 168
rect -19 106 19 142
rect -19 80 -13 106
rect 13 80 19 106
rect -19 44 19 80
rect -19 18 -13 44
rect 13 18 19 44
rect -19 -18 19 18
rect -19 -44 -13 -18
rect 13 -44 19 -18
rect -19 -80 19 -44
rect -19 -106 -13 -80
rect 13 -106 19 -80
rect -19 -142 19 -106
rect -19 -168 -13 -142
rect 13 -168 19 -142
rect -19 -204 19 -168
rect -19 -230 -13 -204
rect 13 -230 19 -204
rect -19 -266 19 -230
rect -19 -292 -13 -266
rect 13 -292 19 -266
rect -19 -328 19 -292
rect -19 -354 -13 -328
rect 13 -354 19 -328
rect -19 -390 19 -354
rect -19 -416 -13 -390
rect 13 -416 19 -390
rect -19 -452 19 -416
rect -19 -478 -13 -452
rect 13 -478 19 -452
rect -19 -514 19 -478
rect -19 -540 -13 -514
rect 13 -540 19 -514
rect -19 -546 19 -540
<< properties >>
string GDS_END 286184
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 284900
<< end >>
