magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 1051 323
<< polysilicon >>
rect -31 182 89 254
rect 193 182 313 254
rect 417 182 537 254
rect 641 182 761 254
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 668 -74 761 -1
use pmos_5p04310590878121_256x8m81  pmos_5p04310590878121_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 1000 302
<< properties >>
string GDS_END 242888
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 242190
<< end >>
