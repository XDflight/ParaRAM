magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -83 3038 3677 6020
rect -83 2098 1171 3038
<< mvnmos >>
rect 3119 1988 3259 2228
rect 335 270 475 1470
rect 579 270 719 1470
rect 823 270 963 1470
rect 1067 270 1207 1470
rect 1311 270 1451 1470
rect 1555 270 1695 1470
rect 1971 270 2111 1470
rect 2215 270 2355 1470
rect 2459 270 2599 1470
rect 2875 270 3015 1470
rect 3119 270 3259 1470
<< mvpmos >>
rect 335 3267 475 5667
rect 579 3267 719 5667
rect 823 3267 963 5667
rect 1067 3267 1207 5667
rect 1483 3267 1623 5667
rect 1727 3267 1867 5667
rect 1971 3267 2111 5667
rect 2387 3267 2527 5667
rect 2631 3267 2771 5667
rect 2875 3267 3015 5667
rect 3119 3267 3259 5667
rect 823 2288 963 2528
<< mvndiff >>
rect 3031 2215 3119 2228
rect 3031 2169 3044 2215
rect 3090 2169 3119 2215
rect 3031 2047 3119 2169
rect 3031 2001 3044 2047
rect 3090 2001 3119 2047
rect 3031 1988 3119 2001
rect 3259 2215 3347 2228
rect 3259 2169 3288 2215
rect 3334 2169 3347 2215
rect 3259 2047 3347 2169
rect 3259 2001 3288 2047
rect 3334 2001 3347 2047
rect 3259 1988 3347 2001
rect 247 1457 335 1470
rect 247 901 260 1457
rect 306 901 335 1457
rect 247 844 335 901
rect 247 798 260 844
rect 306 798 335 844
rect 247 741 335 798
rect 247 695 260 741
rect 306 695 335 741
rect 247 638 335 695
rect 247 592 260 638
rect 306 592 335 638
rect 247 535 335 592
rect 247 489 260 535
rect 306 489 335 535
rect 247 432 335 489
rect 247 386 260 432
rect 306 386 335 432
rect 247 329 335 386
rect 247 283 260 329
rect 306 283 335 329
rect 247 270 335 283
rect 475 1457 579 1470
rect 475 901 504 1457
rect 550 901 579 1457
rect 475 844 579 901
rect 475 798 504 844
rect 550 798 579 844
rect 475 741 579 798
rect 475 695 504 741
rect 550 695 579 741
rect 475 638 579 695
rect 475 592 504 638
rect 550 592 579 638
rect 475 535 579 592
rect 475 489 504 535
rect 550 489 579 535
rect 475 432 579 489
rect 475 386 504 432
rect 550 386 579 432
rect 475 329 579 386
rect 475 283 504 329
rect 550 283 579 329
rect 475 270 579 283
rect 719 1457 823 1470
rect 719 901 748 1457
rect 794 901 823 1457
rect 719 844 823 901
rect 719 798 748 844
rect 794 798 823 844
rect 719 741 823 798
rect 719 695 748 741
rect 794 695 823 741
rect 719 638 823 695
rect 719 592 748 638
rect 794 592 823 638
rect 719 535 823 592
rect 719 489 748 535
rect 794 489 823 535
rect 719 432 823 489
rect 719 386 748 432
rect 794 386 823 432
rect 719 329 823 386
rect 719 283 748 329
rect 794 283 823 329
rect 719 270 823 283
rect 963 1457 1067 1470
rect 963 901 992 1457
rect 1038 901 1067 1457
rect 963 844 1067 901
rect 963 798 992 844
rect 1038 798 1067 844
rect 963 741 1067 798
rect 963 695 992 741
rect 1038 695 1067 741
rect 963 638 1067 695
rect 963 592 992 638
rect 1038 592 1067 638
rect 963 535 1067 592
rect 963 489 992 535
rect 1038 489 1067 535
rect 963 432 1067 489
rect 963 386 992 432
rect 1038 386 1067 432
rect 963 329 1067 386
rect 963 283 992 329
rect 1038 283 1067 329
rect 963 270 1067 283
rect 1207 1457 1311 1470
rect 1207 901 1236 1457
rect 1282 901 1311 1457
rect 1207 844 1311 901
rect 1207 798 1236 844
rect 1282 798 1311 844
rect 1207 741 1311 798
rect 1207 695 1236 741
rect 1282 695 1311 741
rect 1207 638 1311 695
rect 1207 592 1236 638
rect 1282 592 1311 638
rect 1207 535 1311 592
rect 1207 489 1236 535
rect 1282 489 1311 535
rect 1207 432 1311 489
rect 1207 386 1236 432
rect 1282 386 1311 432
rect 1207 329 1311 386
rect 1207 283 1236 329
rect 1282 283 1311 329
rect 1207 270 1311 283
rect 1451 1457 1555 1470
rect 1451 901 1480 1457
rect 1526 901 1555 1457
rect 1451 844 1555 901
rect 1451 798 1480 844
rect 1526 798 1555 844
rect 1451 741 1555 798
rect 1451 695 1480 741
rect 1526 695 1555 741
rect 1451 638 1555 695
rect 1451 592 1480 638
rect 1526 592 1555 638
rect 1451 535 1555 592
rect 1451 489 1480 535
rect 1526 489 1555 535
rect 1451 432 1555 489
rect 1451 386 1480 432
rect 1526 386 1555 432
rect 1451 329 1555 386
rect 1451 283 1480 329
rect 1526 283 1555 329
rect 1451 270 1555 283
rect 1695 1457 1783 1470
rect 1695 901 1724 1457
rect 1770 901 1783 1457
rect 1695 844 1783 901
rect 1695 798 1724 844
rect 1770 798 1783 844
rect 1695 741 1783 798
rect 1695 695 1724 741
rect 1770 695 1783 741
rect 1695 638 1783 695
rect 1695 592 1724 638
rect 1770 592 1783 638
rect 1695 535 1783 592
rect 1695 489 1724 535
rect 1770 489 1783 535
rect 1695 432 1783 489
rect 1695 386 1724 432
rect 1770 386 1783 432
rect 1695 329 1783 386
rect 1695 283 1724 329
rect 1770 283 1783 329
rect 1695 270 1783 283
rect 1883 1457 1971 1470
rect 1883 901 1896 1457
rect 1942 901 1971 1457
rect 1883 844 1971 901
rect 1883 798 1896 844
rect 1942 798 1971 844
rect 1883 741 1971 798
rect 1883 695 1896 741
rect 1942 695 1971 741
rect 1883 638 1971 695
rect 1883 592 1896 638
rect 1942 592 1971 638
rect 1883 535 1971 592
rect 1883 489 1896 535
rect 1942 489 1971 535
rect 1883 432 1971 489
rect 1883 386 1896 432
rect 1942 386 1971 432
rect 1883 329 1971 386
rect 1883 283 1896 329
rect 1942 283 1971 329
rect 1883 270 1971 283
rect 2111 1457 2215 1470
rect 2111 901 2140 1457
rect 2186 901 2215 1457
rect 2111 844 2215 901
rect 2111 798 2140 844
rect 2186 798 2215 844
rect 2111 741 2215 798
rect 2111 695 2140 741
rect 2186 695 2215 741
rect 2111 638 2215 695
rect 2111 592 2140 638
rect 2186 592 2215 638
rect 2111 535 2215 592
rect 2111 489 2140 535
rect 2186 489 2215 535
rect 2111 432 2215 489
rect 2111 386 2140 432
rect 2186 386 2215 432
rect 2111 329 2215 386
rect 2111 283 2140 329
rect 2186 283 2215 329
rect 2111 270 2215 283
rect 2355 1457 2459 1470
rect 2355 901 2384 1457
rect 2430 901 2459 1457
rect 2355 844 2459 901
rect 2355 798 2384 844
rect 2430 798 2459 844
rect 2355 741 2459 798
rect 2355 695 2384 741
rect 2430 695 2459 741
rect 2355 638 2459 695
rect 2355 592 2384 638
rect 2430 592 2459 638
rect 2355 535 2459 592
rect 2355 489 2384 535
rect 2430 489 2459 535
rect 2355 432 2459 489
rect 2355 386 2384 432
rect 2430 386 2459 432
rect 2355 329 2459 386
rect 2355 283 2384 329
rect 2430 283 2459 329
rect 2355 270 2459 283
rect 2599 1457 2687 1470
rect 2599 901 2628 1457
rect 2674 901 2687 1457
rect 2599 844 2687 901
rect 2599 798 2628 844
rect 2674 798 2687 844
rect 2599 741 2687 798
rect 2599 695 2628 741
rect 2674 695 2687 741
rect 2599 638 2687 695
rect 2599 592 2628 638
rect 2674 592 2687 638
rect 2599 535 2687 592
rect 2599 489 2628 535
rect 2674 489 2687 535
rect 2599 432 2687 489
rect 2599 386 2628 432
rect 2674 386 2687 432
rect 2599 329 2687 386
rect 2599 283 2628 329
rect 2674 283 2687 329
rect 2599 270 2687 283
rect 2787 1457 2875 1470
rect 2787 1411 2800 1457
rect 2846 1411 2875 1457
rect 2787 1354 2875 1411
rect 2787 1308 2800 1354
rect 2846 1308 2875 1354
rect 2787 1251 2875 1308
rect 2787 1205 2800 1251
rect 2846 1205 2875 1251
rect 2787 1148 2875 1205
rect 2787 1102 2800 1148
rect 2846 1102 2875 1148
rect 2787 1045 2875 1102
rect 2787 999 2800 1045
rect 2846 999 2875 1045
rect 2787 942 2875 999
rect 2787 896 2800 942
rect 2846 896 2875 942
rect 2787 839 2875 896
rect 2787 283 2800 839
rect 2846 283 2875 839
rect 2787 270 2875 283
rect 3015 1457 3119 1470
rect 3015 1411 3044 1457
rect 3090 1411 3119 1457
rect 3015 1354 3119 1411
rect 3015 1308 3044 1354
rect 3090 1308 3119 1354
rect 3015 1251 3119 1308
rect 3015 1205 3044 1251
rect 3090 1205 3119 1251
rect 3015 1148 3119 1205
rect 3015 1102 3044 1148
rect 3090 1102 3119 1148
rect 3015 1045 3119 1102
rect 3015 999 3044 1045
rect 3090 999 3119 1045
rect 3015 942 3119 999
rect 3015 896 3044 942
rect 3090 896 3119 942
rect 3015 839 3119 896
rect 3015 283 3044 839
rect 3090 283 3119 839
rect 3015 270 3119 283
rect 3259 1457 3347 1470
rect 3259 1411 3288 1457
rect 3334 1411 3347 1457
rect 3259 1354 3347 1411
rect 3259 1308 3288 1354
rect 3334 1308 3347 1354
rect 3259 1251 3347 1308
rect 3259 1205 3288 1251
rect 3334 1205 3347 1251
rect 3259 1148 3347 1205
rect 3259 1102 3288 1148
rect 3334 1102 3347 1148
rect 3259 1045 3347 1102
rect 3259 999 3288 1045
rect 3334 999 3347 1045
rect 3259 942 3347 999
rect 3259 896 3288 942
rect 3334 896 3347 942
rect 3259 839 3347 896
rect 3259 283 3288 839
rect 3334 283 3347 839
rect 3259 270 3347 283
<< mvpdiff >>
rect 247 5654 335 5667
rect 247 3280 260 5654
rect 306 3280 335 5654
rect 247 3267 335 3280
rect 475 5654 579 5667
rect 475 3280 504 5654
rect 550 3280 579 5654
rect 475 3267 579 3280
rect 719 5654 823 5667
rect 719 3280 748 5654
rect 794 3280 823 5654
rect 719 3267 823 3280
rect 963 5654 1067 5667
rect 963 3280 992 5654
rect 1038 3280 1067 5654
rect 963 3267 1067 3280
rect 1207 5654 1295 5667
rect 1207 3280 1236 5654
rect 1282 3280 1295 5654
rect 1207 3267 1295 3280
rect 1395 5654 1483 5667
rect 1395 3280 1408 5654
rect 1454 3280 1483 5654
rect 1395 3267 1483 3280
rect 1623 5654 1727 5667
rect 1623 3280 1652 5654
rect 1698 3280 1727 5654
rect 1623 3267 1727 3280
rect 1867 5654 1971 5667
rect 1867 3280 1896 5654
rect 1942 3280 1971 5654
rect 1867 3267 1971 3280
rect 2111 5654 2199 5667
rect 2111 3280 2140 5654
rect 2186 3280 2199 5654
rect 2111 3267 2199 3280
rect 2299 5654 2387 5667
rect 2299 3280 2312 5654
rect 2358 3280 2387 5654
rect 2299 3267 2387 3280
rect 2527 5654 2631 5667
rect 2527 3280 2556 5654
rect 2602 3280 2631 5654
rect 2527 3267 2631 3280
rect 2771 5654 2875 5667
rect 2771 3280 2800 5654
rect 2846 3280 2875 5654
rect 2771 3267 2875 3280
rect 3015 5654 3119 5667
rect 3015 3280 3044 5654
rect 3090 3280 3119 5654
rect 3015 3267 3119 3280
rect 3259 5654 3347 5667
rect 3259 3280 3288 5654
rect 3334 3280 3347 5654
rect 3259 3267 3347 3280
rect 735 2515 823 2528
rect 735 2469 748 2515
rect 794 2469 823 2515
rect 735 2347 823 2469
rect 735 2301 748 2347
rect 794 2301 823 2347
rect 735 2288 823 2301
rect 963 2515 1051 2528
rect 963 2469 992 2515
rect 1038 2469 1051 2515
rect 963 2347 1051 2469
rect 963 2301 992 2347
rect 1038 2301 1051 2347
rect 963 2288 1051 2301
<< mvndiffc >>
rect 3044 2169 3090 2215
rect 3044 2001 3090 2047
rect 3288 2169 3334 2215
rect 3288 2001 3334 2047
rect 260 901 306 1457
rect 260 798 306 844
rect 260 695 306 741
rect 260 592 306 638
rect 260 489 306 535
rect 260 386 306 432
rect 260 283 306 329
rect 504 901 550 1457
rect 504 798 550 844
rect 504 695 550 741
rect 504 592 550 638
rect 504 489 550 535
rect 504 386 550 432
rect 504 283 550 329
rect 748 901 794 1457
rect 748 798 794 844
rect 748 695 794 741
rect 748 592 794 638
rect 748 489 794 535
rect 748 386 794 432
rect 748 283 794 329
rect 992 901 1038 1457
rect 992 798 1038 844
rect 992 695 1038 741
rect 992 592 1038 638
rect 992 489 1038 535
rect 992 386 1038 432
rect 992 283 1038 329
rect 1236 901 1282 1457
rect 1236 798 1282 844
rect 1236 695 1282 741
rect 1236 592 1282 638
rect 1236 489 1282 535
rect 1236 386 1282 432
rect 1236 283 1282 329
rect 1480 901 1526 1457
rect 1480 798 1526 844
rect 1480 695 1526 741
rect 1480 592 1526 638
rect 1480 489 1526 535
rect 1480 386 1526 432
rect 1480 283 1526 329
rect 1724 901 1770 1457
rect 1724 798 1770 844
rect 1724 695 1770 741
rect 1724 592 1770 638
rect 1724 489 1770 535
rect 1724 386 1770 432
rect 1724 283 1770 329
rect 1896 901 1942 1457
rect 1896 798 1942 844
rect 1896 695 1942 741
rect 1896 592 1942 638
rect 1896 489 1942 535
rect 1896 386 1942 432
rect 1896 283 1942 329
rect 2140 901 2186 1457
rect 2140 798 2186 844
rect 2140 695 2186 741
rect 2140 592 2186 638
rect 2140 489 2186 535
rect 2140 386 2186 432
rect 2140 283 2186 329
rect 2384 901 2430 1457
rect 2384 798 2430 844
rect 2384 695 2430 741
rect 2384 592 2430 638
rect 2384 489 2430 535
rect 2384 386 2430 432
rect 2384 283 2430 329
rect 2628 901 2674 1457
rect 2628 798 2674 844
rect 2628 695 2674 741
rect 2628 592 2674 638
rect 2628 489 2674 535
rect 2628 386 2674 432
rect 2628 283 2674 329
rect 2800 1411 2846 1457
rect 2800 1308 2846 1354
rect 2800 1205 2846 1251
rect 2800 1102 2846 1148
rect 2800 999 2846 1045
rect 2800 896 2846 942
rect 2800 283 2846 839
rect 3044 1411 3090 1457
rect 3044 1308 3090 1354
rect 3044 1205 3090 1251
rect 3044 1102 3090 1148
rect 3044 999 3090 1045
rect 3044 896 3090 942
rect 3044 283 3090 839
rect 3288 1411 3334 1457
rect 3288 1308 3334 1354
rect 3288 1205 3334 1251
rect 3288 1102 3334 1148
rect 3288 999 3334 1045
rect 3288 896 3334 942
rect 3288 283 3334 839
<< mvpdiffc >>
rect 260 3280 306 5654
rect 504 3280 550 5654
rect 748 3280 794 5654
rect 992 3280 1038 5654
rect 1236 3280 1282 5654
rect 1408 3280 1454 5654
rect 1652 3280 1698 5654
rect 1896 3280 1942 5654
rect 2140 3280 2186 5654
rect 2312 3280 2358 5654
rect 2556 3280 2602 5654
rect 2800 3280 2846 5654
rect 3044 3280 3090 5654
rect 3288 3280 3334 5654
rect 748 2469 794 2515
rect 748 2301 794 2347
rect 992 2469 1038 2515
rect 992 2301 1038 2347
<< psubdiff >>
rect 2577 2698 3594 2720
rect 2577 1960 2599 2698
rect 2927 2652 3594 2698
rect 0 1938 2599 1960
rect 2645 2630 3594 2652
rect 0 1892 654 1938
rect 888 1892 2223 1938
rect 2645 1892 2667 2630
rect 3504 2606 3594 2630
rect 0 1870 2667 1892
rect 0 1854 90 1870
rect 0 22 22 1854
rect 68 90 90 1854
rect 3504 90 3526 2606
rect 68 68 3526 90
rect 68 22 176 68
rect 3418 22 3526 68
rect 3572 22 3594 2606
rect 0 0 3594 22
<< nsubdiff >>
rect 0 5915 3594 5937
rect 0 2203 22 5915
rect 68 5869 176 5915
rect 3418 5869 3526 5915
rect 68 5847 3526 5869
rect 68 2203 90 5847
rect 3504 3143 3526 5847
rect 3572 3143 3594 5915
rect 3504 3121 3594 3143
rect 0 2181 90 2203
<< psubdiffcont >>
rect 2599 2652 2927 2698
rect 2599 1938 2645 2652
rect 654 1892 888 1938
rect 2223 1892 2645 1938
rect 22 22 68 1854
rect 176 22 3418 68
rect 3526 22 3572 2606
<< nsubdiffcont >>
rect 22 2203 68 5915
rect 176 5869 3418 5915
rect 3526 3143 3572 5915
<< polysilicon >>
rect 335 5667 475 5711
rect 579 5667 719 5711
rect 823 5667 963 5711
rect 1067 5667 1207 5711
rect 1483 5667 1623 5711
rect 1727 5667 1867 5711
rect 1971 5667 2111 5711
rect 2387 5667 2527 5711
rect 2631 5667 2771 5711
rect 2875 5667 3015 5711
rect 3119 5667 3259 5711
rect 335 3089 475 3267
rect 579 3089 719 3267
rect 335 3070 719 3089
rect 335 3024 416 3070
rect 650 3024 719 3070
rect 335 3005 719 3024
rect 823 3089 963 3267
rect 1067 3089 1207 3267
rect 823 3070 1207 3089
rect 823 3024 906 3070
rect 1140 3024 1207 3070
rect 823 3005 1207 3024
rect 1483 3070 1623 3267
rect 1483 2930 1530 3070
rect 1576 2930 1623 3070
rect 1483 2911 1623 2930
rect 1727 3070 1867 3267
rect 1727 2930 1774 3070
rect 1820 2930 1867 3070
rect 1727 2911 1867 2930
rect 1971 3070 2111 3267
rect 2387 3207 2527 3267
rect 2631 3207 2771 3267
rect 2875 3207 3015 3267
rect 3119 3207 3259 3267
rect 2387 3188 3259 3207
rect 2387 3142 2706 3188
rect 2940 3142 3259 3188
rect 2387 3123 3259 3142
rect 1971 2930 2018 3070
rect 2064 2930 2111 3070
rect 1971 2911 2111 2930
rect 823 2528 963 2572
rect 823 2228 963 2288
rect 757 2209 963 2228
rect 757 2163 776 2209
rect 916 2163 963 2209
rect 757 2144 963 2163
rect 3119 2431 3259 2450
rect 3119 2291 3166 2431
rect 3212 2291 3259 2431
rect 3119 2228 3259 2291
rect 3119 1944 3259 1988
rect 335 1673 1207 1692
rect 335 1533 382 1673
rect 428 1533 1114 1673
rect 1160 1533 1207 1673
rect 335 1530 1207 1533
rect 335 1470 475 1530
rect 579 1470 719 1530
rect 823 1470 963 1530
rect 1067 1470 1207 1530
rect 1311 1673 1451 1692
rect 1311 1533 1358 1673
rect 1404 1533 1451 1673
rect 1311 1470 1451 1533
rect 1555 1673 1695 1692
rect 1555 1533 1602 1673
rect 1648 1533 1695 1673
rect 1555 1470 1695 1533
rect 1971 1673 2111 1692
rect 1971 1533 2018 1673
rect 2064 1533 2111 1673
rect 1971 1470 2111 1533
rect 2215 1673 2599 1692
rect 2215 1533 2262 1673
rect 2308 1533 2599 1673
rect 2215 1530 2599 1533
rect 2215 1470 2355 1530
rect 2459 1470 2599 1530
rect 2875 1673 3259 1692
rect 2875 1533 2922 1673
rect 2968 1533 3259 1673
rect 2875 1530 3259 1533
rect 2875 1470 3015 1530
rect 3119 1470 3259 1530
rect 335 226 475 270
rect 579 226 719 270
rect 823 226 963 270
rect 1067 226 1207 270
rect 1311 226 1451 270
rect 1555 226 1695 270
rect 1971 226 2111 270
rect 2215 226 2355 270
rect 2459 226 2599 270
rect 2875 226 3015 270
rect 3119 226 3259 270
<< polycontact >>
rect 416 3024 650 3070
rect 906 3024 1140 3070
rect 1530 2930 1576 3070
rect 1774 2930 1820 3070
rect 2706 3142 2940 3188
rect 2018 2930 2064 3070
rect 776 2163 916 2209
rect 3166 2291 3212 2431
rect 382 1533 428 1673
rect 1114 1533 1160 1673
rect 1358 1533 1404 1673
rect 1602 1533 1648 1673
rect 2018 1533 2064 1673
rect 2262 1533 2308 1673
rect 2922 1533 2968 1673
<< metal1 >>
rect 11 5915 3583 5926
rect 11 2203 22 5915
rect 68 5869 176 5915
rect 3418 5869 3526 5915
rect 68 5858 3526 5869
rect 68 2203 79 5858
rect 245 5654 321 5667
rect 245 3280 260 5654
rect 306 3280 321 5654
rect 245 3217 321 3280
rect 489 5654 565 5858
rect 489 3280 504 5654
rect 550 3280 565 5654
rect 489 3267 565 3280
rect 733 5654 809 5667
rect 733 3280 748 5654
rect 794 3280 809 5654
rect 733 3217 809 3280
rect 977 5654 1053 5667
rect 977 3435 992 5654
rect 1038 3435 1053 5654
rect 977 3279 989 3435
rect 1041 3279 1053 3435
rect 977 3267 1053 3279
rect 1221 5654 1297 5667
rect 1221 3280 1236 5654
rect 1282 3280 1297 5654
rect 1221 3217 1297 3280
rect 245 3141 1297 3217
rect 11 2192 79 2203
rect 367 3070 661 3081
rect 367 3024 416 3070
rect 650 3024 661 3070
rect 367 3013 661 3024
rect 831 3070 1151 3081
rect 831 3069 906 3070
rect 11 1854 79 1865
rect 11 22 22 1854
rect 68 79 79 1854
rect 367 1673 443 3013
rect 831 2913 843 3069
rect 895 3024 906 3069
rect 1140 3024 1151 3070
rect 895 3013 1151 3024
rect 895 2913 907 3013
rect 831 2901 907 2913
rect 977 2881 1053 2893
rect 977 2789 989 2881
rect 367 1533 382 1673
rect 428 1533 443 1673
rect 367 1522 443 1533
rect 489 2725 989 2789
rect 1041 2725 1053 2881
rect 489 2713 1053 2725
rect 489 2528 565 2713
rect 1221 2528 1297 3141
rect 1393 5654 1469 5667
rect 1393 3280 1408 5654
rect 1454 3280 1469 5654
rect 1393 3173 1469 3280
rect 1393 3017 1405 3173
rect 1457 3017 1469 3173
rect 1637 5654 1713 5667
rect 1637 3280 1652 5654
rect 1698 3280 1713 5654
rect 1637 3217 1713 3280
rect 1881 5654 1957 5858
rect 1881 3280 1896 5654
rect 1942 3280 1957 5654
rect 1881 3267 1957 3280
rect 2125 5654 2201 5667
rect 2125 3280 2140 5654
rect 2186 3280 2201 5654
rect 2125 3217 2201 3280
rect 2297 5654 2373 5858
rect 2297 3280 2312 5654
rect 2358 3280 2373 5654
rect 2297 3267 2373 3280
rect 2529 5654 2629 5667
rect 2529 3280 2556 5654
rect 2602 3280 2629 5654
rect 1637 3141 2201 3217
rect 1393 3005 1469 3017
rect 1515 3070 1591 3081
rect 1515 2930 1530 3070
rect 1576 2930 1591 3070
rect 1515 2652 1591 2930
rect 489 2515 794 2528
rect 489 2469 748 2515
rect 489 2347 794 2469
rect 489 2301 748 2347
rect 489 2288 794 2301
rect 977 2515 1297 2528
rect 977 2469 992 2515
rect 1038 2469 1297 2515
rect 977 2452 1297 2469
rect 1343 2576 1591 2652
rect 1637 3069 1713 3081
rect 1637 2913 1649 3069
rect 1701 2913 1713 3069
rect 977 2347 1053 2452
rect 977 2301 992 2347
rect 1038 2301 1053 2347
rect 245 1457 321 1470
rect 245 901 260 1457
rect 306 901 321 1457
rect 245 844 321 901
rect 245 798 260 844
rect 306 798 321 844
rect 245 741 321 798
rect 245 695 260 741
rect 306 695 321 741
rect 245 638 321 695
rect 245 592 260 638
rect 306 592 321 638
rect 245 535 321 592
rect 245 489 260 535
rect 306 489 321 535
rect 245 432 321 489
rect 245 386 260 432
rect 306 386 321 432
rect 245 329 321 386
rect 245 283 260 329
rect 306 283 321 329
rect 245 79 321 283
rect 489 1457 565 2288
rect 733 2209 927 2220
rect 733 2163 776 2209
rect 916 2163 927 2209
rect 733 2152 927 2163
rect 733 1949 809 2152
rect 643 1938 899 1949
rect 643 1892 654 1938
rect 888 1892 899 1938
rect 643 1881 899 1892
rect 489 901 504 1457
rect 550 901 565 1457
rect 489 844 565 901
rect 489 798 504 844
rect 550 798 565 844
rect 489 741 565 798
rect 489 695 504 741
rect 550 695 565 741
rect 489 638 565 695
rect 489 592 504 638
rect 550 592 565 638
rect 489 535 565 592
rect 489 489 504 535
rect 550 489 565 535
rect 489 432 565 489
rect 489 386 504 432
rect 550 386 565 432
rect 489 329 565 386
rect 489 283 504 329
rect 550 283 565 329
rect 489 270 565 283
rect 733 1457 809 1881
rect 733 901 748 1457
rect 794 901 809 1457
rect 733 844 809 901
rect 733 798 748 844
rect 794 798 809 844
rect 733 741 809 798
rect 733 695 748 741
rect 794 695 809 741
rect 733 638 809 695
rect 733 592 748 638
rect 794 592 809 638
rect 733 535 809 592
rect 733 489 748 535
rect 794 489 809 535
rect 733 432 809 489
rect 733 386 748 432
rect 794 386 809 432
rect 733 329 809 386
rect 733 283 748 329
rect 794 283 809 329
rect 733 79 809 283
rect 977 1457 1053 2301
rect 1099 2202 1175 2214
rect 1099 2046 1111 2202
rect 1163 2046 1175 2202
rect 1099 1673 1175 2046
rect 1099 1533 1114 1673
rect 1160 1533 1175 1673
rect 1099 1522 1175 1533
rect 1343 1673 1419 2576
rect 1637 2494 1713 2913
rect 1343 1533 1358 1673
rect 1404 1533 1419 1673
rect 1343 1522 1419 1533
rect 1465 2418 1713 2494
rect 1759 3070 1835 3081
rect 1759 2930 1774 3070
rect 1820 2930 1835 3070
rect 977 901 992 1457
rect 1038 901 1053 1457
rect 977 844 1053 901
rect 977 798 992 844
rect 1038 798 1053 844
rect 977 741 1053 798
rect 977 695 992 741
rect 1038 695 1053 741
rect 977 638 1053 695
rect 977 592 992 638
rect 1038 592 1053 638
rect 977 535 1053 592
rect 977 489 992 535
rect 1038 489 1053 535
rect 977 432 1053 489
rect 977 386 992 432
rect 1038 386 1053 432
rect 977 329 1053 386
rect 977 283 992 329
rect 1038 283 1053 329
rect 977 270 1053 283
rect 1221 1457 1297 1470
rect 1221 901 1236 1457
rect 1282 901 1297 1457
rect 1221 844 1297 901
rect 1221 798 1236 844
rect 1282 798 1297 844
rect 1221 741 1297 798
rect 1221 695 1236 741
rect 1282 695 1297 741
rect 1221 638 1297 695
rect 1221 592 1236 638
rect 1282 592 1297 638
rect 1221 535 1297 592
rect 1221 489 1236 535
rect 1282 489 1297 535
rect 1221 432 1297 489
rect 1221 386 1236 432
rect 1282 386 1297 432
rect 1221 329 1297 386
rect 1221 283 1236 329
rect 1282 283 1297 329
rect 1221 79 1297 283
rect 1465 1457 1541 2418
rect 1759 2350 1835 2930
rect 1587 2274 1835 2350
rect 1587 1673 1663 2274
rect 1881 2110 1957 3141
rect 1587 1533 1602 1673
rect 1648 1533 1663 1673
rect 1587 1522 1663 1533
rect 1709 2098 1957 2110
rect 1709 2046 1755 2098
rect 1911 2046 1957 2098
rect 1709 2034 1957 2046
rect 2003 3070 2079 3081
rect 2003 2930 2018 3070
rect 2064 2930 2079 3070
rect 1465 901 1480 1457
rect 1526 901 1541 1457
rect 1465 844 1541 901
rect 1465 798 1480 844
rect 1526 798 1541 844
rect 1465 741 1541 798
rect 1465 695 1480 741
rect 1526 695 1541 741
rect 1465 638 1541 695
rect 1465 592 1480 638
rect 1526 592 1541 638
rect 1465 535 1541 592
rect 1465 489 1480 535
rect 1526 489 1541 535
rect 1465 432 1541 489
rect 1465 386 1480 432
rect 1526 386 1541 432
rect 1465 329 1541 386
rect 1465 283 1480 329
rect 1526 283 1541 329
rect 1465 212 1541 283
rect 1709 1457 1785 2034
rect 2003 1673 2079 2930
rect 2529 2945 2629 3280
rect 2785 5654 2861 5858
rect 2785 3280 2800 5654
rect 2846 3280 2861 5654
rect 2785 3267 2861 3280
rect 3017 5654 3117 5667
rect 3017 3280 3044 5654
rect 3090 3280 3117 5654
rect 2695 3188 2951 3199
rect 2695 3142 2706 3188
rect 2940 3142 2951 3188
rect 2695 3069 2951 3142
rect 2695 3017 2745 3069
rect 2901 3017 2951 3069
rect 2695 3005 2951 3017
rect 3017 3105 3117 3280
rect 3273 5654 3349 5858
rect 3273 3485 3288 5654
rect 3334 3485 3349 5654
rect 3273 3329 3285 3485
rect 3337 3329 3349 3485
rect 3273 3280 3288 3329
rect 3334 3280 3349 3329
rect 3273 3267 3349 3280
rect 3515 3143 3526 5858
rect 3572 3143 3583 5915
rect 3515 3132 3583 3143
rect 3017 3005 3373 3105
rect 2529 2845 3105 2945
rect 2588 2698 2938 2709
rect 2588 1953 2599 2698
rect 2927 2652 2938 2698
rect 2003 1533 2018 1673
rect 2064 1533 2079 1673
rect 2003 1522 2079 1533
rect 2125 1941 2599 1953
rect 2645 2641 2938 2652
rect 2125 1938 2280 1941
rect 2125 1892 2223 1938
rect 2645 1892 2656 2641
rect 2125 1889 2280 1892
rect 2644 1889 2656 1892
rect 2125 1877 2656 1889
rect 3029 2215 3105 2845
rect 3151 2448 3227 2460
rect 3151 2292 3163 2448
rect 3215 2292 3227 2448
rect 3151 2291 3166 2292
rect 3212 2291 3227 2292
rect 3151 2280 3227 2291
rect 3029 2169 3044 2215
rect 3090 2169 3105 2215
rect 3029 2047 3105 2169
rect 3029 2001 3044 2047
rect 3090 2001 3105 2047
rect 1709 901 1724 1457
rect 1770 901 1785 1457
rect 1709 844 1785 901
rect 1709 798 1724 844
rect 1770 798 1785 844
rect 1709 741 1785 798
rect 1709 695 1724 741
rect 1770 695 1785 741
rect 1709 638 1785 695
rect 1709 592 1724 638
rect 1770 592 1785 638
rect 1709 535 1785 592
rect 1709 489 1724 535
rect 1770 489 1785 535
rect 1709 432 1785 489
rect 1709 386 1724 432
rect 1770 386 1785 432
rect 1709 329 1785 386
rect 1709 283 1724 329
rect 1770 283 1785 329
rect 1709 270 1785 283
rect 1881 1457 1957 1470
rect 1881 901 1896 1457
rect 1942 901 1957 1457
rect 1881 844 1957 901
rect 1881 798 1896 844
rect 1942 798 1957 844
rect 1881 741 1957 798
rect 1881 695 1896 741
rect 1942 695 1957 741
rect 1881 638 1957 695
rect 1881 592 1896 638
rect 1942 592 1957 638
rect 1881 535 1957 592
rect 1881 489 1896 535
rect 1942 489 1957 535
rect 1881 432 1957 489
rect 1881 386 1896 432
rect 1942 386 1957 432
rect 1881 329 1957 386
rect 1881 283 1896 329
rect 1942 283 1957 329
rect 1881 212 1957 283
rect 2125 1457 2201 1877
rect 3029 1824 3105 2001
rect 2369 1748 3105 1824
rect 2125 901 2140 1457
rect 2186 901 2201 1457
rect 2125 844 2201 901
rect 2125 798 2140 844
rect 2186 798 2201 844
rect 2125 741 2201 798
rect 2125 695 2140 741
rect 2186 695 2201 741
rect 2125 638 2201 695
rect 2125 592 2140 638
rect 2186 592 2201 638
rect 2125 535 2201 592
rect 2125 489 2140 535
rect 2186 489 2201 535
rect 2125 432 2201 489
rect 2125 386 2140 432
rect 2186 386 2201 432
rect 2125 329 2201 386
rect 2125 283 2140 329
rect 2186 283 2201 329
rect 2125 270 2201 283
rect 2247 1673 2323 1684
rect 2247 1533 2262 1673
rect 2308 1533 2323 1673
rect 2247 212 2323 1533
rect 2369 1457 2445 1748
rect 2907 1690 2983 1702
rect 2907 1534 2919 1690
rect 2971 1534 2983 1690
rect 2907 1533 2922 1534
rect 2968 1533 2983 1534
rect 2907 1522 2983 1533
rect 2369 901 2384 1457
rect 2430 901 2445 1457
rect 2369 844 2445 901
rect 2369 798 2384 844
rect 2430 798 2445 844
rect 2369 741 2445 798
rect 2369 695 2384 741
rect 2430 695 2445 741
rect 2369 638 2445 695
rect 2369 592 2384 638
rect 2430 592 2445 638
rect 2369 535 2445 592
rect 2369 489 2384 535
rect 2430 489 2445 535
rect 2369 432 2445 489
rect 2369 386 2384 432
rect 2430 386 2445 432
rect 2369 329 2445 386
rect 2369 283 2384 329
rect 2430 283 2445 329
rect 2369 270 2445 283
rect 2613 1457 2689 1470
rect 2613 901 2628 1457
rect 2674 901 2689 1457
rect 2613 844 2689 901
rect 2613 798 2628 844
rect 2674 798 2689 844
rect 2613 741 2689 798
rect 2613 695 2628 741
rect 2674 695 2689 741
rect 2613 638 2689 695
rect 2613 592 2628 638
rect 2674 592 2689 638
rect 2613 535 2689 592
rect 2613 489 2628 535
rect 2674 489 2689 535
rect 2613 432 2689 489
rect 2613 386 2628 432
rect 2674 386 2689 432
rect 2613 329 2689 386
rect 2613 283 2628 329
rect 2674 283 2689 329
rect 1465 136 2323 212
rect 2613 79 2689 283
rect 2773 1457 2873 1470
rect 2773 1411 2800 1457
rect 2846 1411 2873 1457
rect 2773 1354 2873 1411
rect 2773 1308 2800 1354
rect 2846 1308 2873 1354
rect 2773 1251 2873 1308
rect 2773 1205 2800 1251
rect 2846 1205 2873 1251
rect 2773 1148 2873 1205
rect 2773 1102 2800 1148
rect 2846 1102 2873 1148
rect 2773 1045 2873 1102
rect 2773 999 2800 1045
rect 2846 999 2873 1045
rect 2773 942 2873 999
rect 2773 896 2800 942
rect 2846 896 2873 942
rect 2773 839 2873 896
rect 2773 283 2800 839
rect 2846 283 2873 839
rect 2773 219 2873 283
rect 3029 1457 3105 1748
rect 3029 1411 3044 1457
rect 3090 1411 3105 1457
rect 3029 1354 3105 1411
rect 3029 1308 3044 1354
rect 3090 1308 3105 1354
rect 3029 1251 3105 1308
rect 3029 1205 3044 1251
rect 3090 1205 3105 1251
rect 3029 1148 3105 1205
rect 3029 1102 3044 1148
rect 3090 1102 3105 1148
rect 3029 1045 3105 1102
rect 3029 999 3044 1045
rect 3090 999 3105 1045
rect 3029 942 3105 999
rect 3029 896 3044 942
rect 3090 896 3105 942
rect 3029 839 3105 896
rect 3029 283 3044 839
rect 3090 283 3105 839
rect 3029 270 3105 283
rect 3273 2215 3373 3005
rect 3445 2641 3583 2709
rect 3273 2169 3288 2215
rect 3334 2169 3373 2215
rect 3273 2047 3373 2169
rect 3273 2001 3288 2047
rect 3334 2001 3373 2047
rect 3273 1457 3373 2001
rect 3273 1411 3288 1457
rect 3334 1411 3373 1457
rect 3273 1354 3373 1411
rect 3273 1308 3288 1354
rect 3334 1308 3373 1354
rect 3273 1251 3373 1308
rect 3273 1205 3288 1251
rect 3334 1205 3373 1251
rect 3273 1148 3373 1205
rect 3273 1102 3288 1148
rect 3334 1102 3373 1148
rect 3273 1045 3373 1102
rect 3273 999 3288 1045
rect 3334 999 3373 1045
rect 3273 942 3373 999
rect 3273 896 3288 942
rect 3334 896 3373 942
rect 3273 839 3373 896
rect 3273 283 3288 839
rect 3334 283 3373 839
rect 3273 219 3373 283
rect 2773 129 3373 219
rect 3515 2606 3583 2641
rect 3515 79 3526 2606
rect 68 68 3526 79
rect 68 22 176 68
rect 3418 22 3526 68
rect 3572 22 3583 2606
rect 11 11 3583 22
<< via1 >>
rect 989 3280 992 3435
rect 992 3280 1038 3435
rect 1038 3280 1041 3435
rect 989 3279 1041 3280
rect 843 2913 895 3069
rect 989 2725 1041 2881
rect 1405 3017 1457 3173
rect 1649 2913 1701 3069
rect 1111 2046 1163 2202
rect 1755 2046 1911 2098
rect 2745 3017 2901 3069
rect 3285 3329 3288 3485
rect 3288 3329 3334 3485
rect 3334 3329 3337 3485
rect 2280 1938 2599 1941
rect 2599 1938 2644 1941
rect 2280 1892 2644 1938
rect 2280 1889 2644 1892
rect 3163 2431 3215 2448
rect 3163 2292 3166 2431
rect 3166 2292 3212 2431
rect 3212 2292 3215 2431
rect 2919 1673 2971 1690
rect 2919 1534 2922 1673
rect 2922 1534 2968 1673
rect 2968 1534 2971 1673
<< metal2 >>
rect 3273 3485 3349 3497
rect 977 3435 1053 3447
rect 977 3279 989 3435
rect 1041 3279 1053 3435
rect 831 3069 907 3081
rect 831 2913 843 3069
rect 895 2913 907 3069
rect 831 2901 907 2913
rect 977 2881 1053 3279
rect 3273 3329 3285 3485
rect 3337 3329 3349 3485
rect 1393 3173 1469 3185
rect 1393 3017 1405 3173
rect 1457 3081 1469 3173
rect 1457 3069 2951 3081
rect 1457 3017 1649 3069
rect 1393 3005 1649 3017
rect 1637 2913 1649 3005
rect 1701 3017 2745 3069
rect 2901 3017 2951 3069
rect 1701 3005 2951 3017
rect 1701 2913 1713 3005
rect 1637 2901 1713 2913
rect 977 2725 989 2881
rect 1041 2725 1053 2881
rect 977 2713 1053 2725
rect 3273 2460 3349 3329
rect 3151 2448 3349 2460
rect 3151 2292 3163 2448
rect 3215 2292 3349 2448
rect 3151 2280 3349 2292
rect 1099 2202 1175 2214
rect 1099 2046 1111 2202
rect 1163 2110 1175 2202
rect 1163 2098 1957 2110
rect 1163 2046 1755 2098
rect 1911 2046 1957 2098
rect 1099 2034 1957 2046
rect 2268 1941 3549 1953
rect 2268 1889 2280 1941
rect 2644 1889 3549 1941
rect 2268 1877 3549 1889
rect 2907 1690 2983 1702
rect 2907 1534 2919 1690
rect 2971 1534 2983 1690
rect 2907 1522 2983 1534
use M1_NWELL_CDNS_40661954729417  M1_NWELL_CDNS_40661954729417_0
timestamp 1666464484
transform 1 0 3549 0 1 4529
box 0 0 1 1
use M1_NWELL_CDNS_40661954729472  M1_NWELL_CDNS_40661954729472_0
timestamp 1666464484
transform 1 0 1797 0 1 5892
box 0 0 1 1
use M1_NWELL_CDNS_40661954729477  M1_NWELL_CDNS_40661954729477_0
timestamp 1666464484
transform 1 0 45 0 1 4059
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_0
timestamp 1666464484
transform 0 -1 1797 -1 0 3000
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_1
timestamp 1666464484
transform 0 -1 2041 -1 0 3000
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_2
timestamp 1666464484
transform 0 -1 1553 -1 0 3000
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_3
timestamp 1666464484
transform 0 -1 2041 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_4
timestamp 1666464484
transform 0 -1 2945 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_5
timestamp 1666464484
transform 0 -1 2285 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_6
timestamp 1666464484
transform 0 -1 1381 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_7
timestamp 1666464484
transform 0 -1 1137 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_8
timestamp 1666464484
transform 0 -1 1625 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_9
timestamp 1666464484
transform 0 -1 3189 1 0 2361
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_10
timestamp 1666464484
transform 0 -1 405 1 0 1603
box 0 0 1 1
use M1_POLY2_CDNS_40661954729255  M1_POLY2_CDNS_40661954729255_11
timestamp 1666464484
transform 1 0 846 0 1 2186
box 0 0 1 1
use M1_POLY2_CDNS_40661954729471  M1_POLY2_CDNS_40661954729471_0
timestamp 1666464484
transform 1 0 533 0 -1 3047
box 0 0 1 1
use M1_POLY2_CDNS_40661954729471  M1_POLY2_CDNS_40661954729471_1
timestamp 1666464484
transform 1 0 1023 0 -1 3047
box 0 0 1 1
use M1_POLY2_CDNS_40661954729471  M1_POLY2_CDNS_40661954729471_2
timestamp 1666464484
transform -1 0 2823 0 -1 3165
box 0 0 1 1
use M1_PSUB_CDNS_40661954729416  M1_PSUB_CDNS_40661954729416_0
timestamp 1666464484
transform 1 0 2434 0 1 1915
box 0 0 1 1
use M1_PSUB_CDNS_40661954729473  M1_PSUB_CDNS_40661954729473_0
timestamp 1666464484
transform 1 0 1797 0 1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661954729474  M1_PSUB_CDNS_40661954729474_0
timestamp 1666464484
transform 1 0 2763 0 1 2675
box 0 0 1 1
use M1_PSUB_CDNS_40661954729475  M1_PSUB_CDNS_40661954729475_0
timestamp 1666464484
transform 1 0 3549 0 1 1314
box 0 0 1 1
use M1_PSUB_CDNS_40661954729476  M1_PSUB_CDNS_40661954729476_0
timestamp 1666464484
transform 1 0 771 0 1 1915
box 0 0 1 1
use M1_PSUB_CDNS_40661954729478  M1_PSUB_CDNS_40661954729478_0
timestamp 1666464484
transform 1 0 2622 0 1 2297
box 0 0 1 1
use M1_PSUB_CDNS_40661954729479  M1_PSUB_CDNS_40661954729479_0
timestamp 1666464484
transform 1 0 45 0 1 938
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_0
timestamp 1666464484
transform 0 -1 2823 1 0 3043
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_1
timestamp 1666464484
transform 0 -1 1833 1 0 2072
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_2
timestamp 1666464484
transform 1 0 1137 0 1 2124
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_3
timestamp 1666464484
transform 1 0 1015 0 1 2803
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_4
timestamp 1666464484
transform 1 0 3311 0 1 3407
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_5
timestamp 1666464484
transform 1 0 3189 0 1 2370
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_6
timestamp 1666464484
transform 1 0 2945 0 1 1612
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_7
timestamp 1666464484
transform 1 0 1431 0 1 3095
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_8
timestamp 1666464484
transform 1 0 1015 0 1 3357
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_9
timestamp 1666464484
transform 1 0 869 0 1 2991
box 0 0 1 1
use M2_M1_CDNS_40661954729341  M2_M1_CDNS_40661954729341_10
timestamp 1666464484
transform 1 0 1675 0 1 2991
box 0 0 1 1
use M2_M1_CDNS_40661954729407  M2_M1_CDNS_40661954729407_0
timestamp 1666464484
transform 1 0 2462 0 1 1915
box 0 0 1 1
use nmos_6p0_CDNS_4066195472940  nmos_6p0_CDNS_4066195472940_0
timestamp 1666464484
transform 1 0 3119 0 1 1988
box 0 0 1 1
use nmos_6p0_CDNS_4066195472944  nmos_6p0_CDNS_4066195472944_0
timestamp 1666464484
transform -1 0 1207 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472944  nmos_6p0_CDNS_4066195472944_1
timestamp 1666464484
transform -1 0 2599 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472945  nmos_6p0_CDNS_4066195472945_0
timestamp 1666464484
transform -1 0 2111 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472945  nmos_6p0_CDNS_4066195472945_1
timestamp 1666464484
transform -1 0 1451 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472945  nmos_6p0_CDNS_4066195472945_2
timestamp 1666464484
transform -1 0 1695 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472946  nmos_6p0_CDNS_4066195472946_0
timestamp 1666464484
transform -1 0 719 0 1 270
box 0 0 1 1
use nmos_6p0_CDNS_4066195472946  nmos_6p0_CDNS_4066195472946_1
timestamp 1666464484
transform -1 0 3259 0 -1 1470
box 0 0 1 1
use pmos_6p0_CDNS_4066195472941  pmos_6p0_CDNS_4066195472941_0
timestamp 1666464484
transform -1 0 2111 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472941  pmos_6p0_CDNS_4066195472941_1
timestamp 1666464484
transform -1 0 1623 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472941  pmos_6p0_CDNS_4066195472941_2
timestamp 1666464484
transform -1 0 1867 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472942  pmos_6p0_CDNS_4066195472942_0
timestamp 1666464484
transform 1 0 335 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472942  pmos_6p0_CDNS_4066195472942_1
timestamp 1666464484
transform 1 0 2875 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472942  pmos_6p0_CDNS_4066195472942_2
timestamp 1666464484
transform 1 0 2387 0 1 3267
box 0 0 1 1
use pmos_6p0_CDNS_4066195472943  pmos_6p0_CDNS_4066195472943_0
timestamp 1666464484
transform -1 0 963 0 1 2288
box 0 0 1 1
use pmos_6p0_CDNS_4066195472947  pmos_6p0_CDNS_4066195472947_0
timestamp 1666464484
transform -1 0 1207 0 -1 5667
box 0 0 1 1
<< labels >>
rlabel metal2 s 869 3046 869 3046 4 SL
port 1 nsew
rlabel metal2 s 2947 1602 2947 1602 4 SLB
port 2 nsew
rlabel metal1 s 1015 5270 1015 5270 4 NDRIVE_X
port 3 nsew
rlabel metal1 s 1390 1726 1390 1726 4 ENB
port 4 nsew
rlabel metal1 s 284 47 284 47 4 DVSS
port 5 nsew
rlabel metal1 s 2042 1726 2042 1726 4 A
port 6 nsew
rlabel metal1 s 345 5891 345 5891 4 DVDD
port 7 nsew
rlabel metal1 s 772 5265 772 5265 4 NDRIVE_Y
port 8 nsew
rlabel metal1 s 2580 5278 2580 5278 4 PDRIVE_Y
port 9 nsew
rlabel metal1 s 3066 5296 3066 5296 4 PDRIVE_X
port 10 nsew
rlabel metal1 s 1632 1726 1632 1726 4 EN
port 11 nsew
<< properties >>
string GDS_END 1854340
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1844998
string path 25.375 86.175 25.375 67.825 
<< end >>
