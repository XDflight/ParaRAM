magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 2464 844
rect 273 610 319 724
rect 354 424 430 550
rect 165 360 430 424
rect 697 617 743 724
rect 273 60 319 163
rect 670 248 886 312
rect 677 60 723 165
rect 800 110 886 248
rect 1482 561 1550 724
rect 1941 506 1987 724
rect 1553 60 1599 179
rect 1921 60 1967 211
rect 2132 106 2216 676
rect 2349 506 2395 724
rect 2369 60 2415 211
rect 0 -60 2464 60
<< obsm1 >>
rect 38 278 115 678
rect 522 417 579 678
rect 1020 628 1301 674
rect 625 467 1020 513
rect 1151 417 1197 562
rect 522 371 1197 417
rect 38 232 472 278
rect 38 106 115 232
rect 522 106 590 371
rect 957 202 1003 371
rect 1255 295 1301 628
rect 1697 461 1743 645
rect 1364 415 1834 461
rect 1255 249 1716 295
rect 1255 152 1301 249
rect 1040 106 1301 152
rect 1766 106 1834 415
<< labels >>
rlabel metal1 s 670 248 886 312 6 D
port 1 nsew default input
rlabel metal1 s 800 110 886 248 6 D
port 1 nsew default input
rlabel metal1 s 354 424 430 550 6 E
port 2 nsew clock input
rlabel metal1 s 165 360 430 424 6 E
port 2 nsew clock input
rlabel metal1 s 2132 106 2216 676 6 Q
port 3 nsew default output
rlabel metal1 s 0 724 2464 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 617 2395 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 617 1987 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 617 1550 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 697 617 743 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 617 319 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 610 2395 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 610 1987 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 610 1550 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 610 319 617 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 561 2395 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 561 1987 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1482 561 1550 610 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2349 506 2395 561 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1941 506 1987 561 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2369 179 2415 211 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 179 1967 211 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 165 2415 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 165 1967 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 165 1599 179 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 163 2415 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 163 1967 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 163 1599 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 163 723 165 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2369 60 2415 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1921 60 1967 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1553 60 1599 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 677 60 723 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 163 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2464 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 580594
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 574928
<< end >>
