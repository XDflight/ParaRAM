magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -170 681 170 716
rect -170 625 -134 681
rect -78 625 78 681
rect 134 625 170 681
rect -170 463 170 625
rect -170 407 -134 463
rect -78 407 78 463
rect 134 407 170 463
rect -170 246 170 407
rect -170 190 -134 246
rect -78 190 78 246
rect 134 190 170 246
rect -170 28 170 190
rect -170 -28 -134 28
rect -78 -28 78 28
rect 134 -28 170 28
rect -170 -190 170 -28
rect -170 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 170 -190
rect -170 -407 170 -246
rect -170 -463 -134 -407
rect -78 -463 78 -407
rect 134 -463 170 -407
rect -170 -625 170 -463
rect -170 -681 -134 -625
rect -78 -681 78 -625
rect 134 -681 170 -625
rect -170 -843 170 -681
rect -170 -899 -134 -843
rect -78 -899 78 -843
rect 134 -899 170 -843
rect -170 -1060 170 -899
rect -170 -1116 -134 -1060
rect -78 -1116 78 -1060
rect 134 -1116 170 -1060
rect -170 -1155 170 -1116
<< via2 >>
rect -134 625 -78 681
rect 78 625 134 681
rect -134 407 -78 463
rect 78 407 134 463
rect -134 190 -78 246
rect 78 190 134 246
rect -134 -28 -78 28
rect 78 -28 134 28
rect -134 -246 -78 -190
rect 78 -246 134 -190
rect -134 -463 -78 -407
rect 78 -463 134 -407
rect -134 -681 -78 -625
rect 78 -681 134 -625
rect -134 -899 -78 -843
rect 78 -899 134 -843
rect -134 -1116 -78 -1060
rect 78 -1116 134 -1060
<< metal3 >>
rect -170 681 170 716
rect -170 625 -134 681
rect -78 625 78 681
rect 134 625 170 681
rect -170 463 170 625
rect -170 407 -134 463
rect -78 407 78 463
rect 134 407 170 463
rect -170 246 170 407
rect -170 190 -134 246
rect -78 190 78 246
rect 134 190 170 246
rect -170 28 170 190
rect -170 -28 -134 28
rect -78 -28 78 28
rect 134 -28 170 28
rect -170 -190 170 -28
rect -170 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 170 -190
rect -170 -407 170 -246
rect -170 -463 -134 -407
rect -78 -463 78 -407
rect 134 -463 170 -407
rect -170 -625 170 -463
rect -170 -681 -134 -625
rect -78 -681 78 -625
rect 134 -681 170 -625
rect -170 -843 170 -681
rect -170 -899 -134 -843
rect -78 -899 78 -843
rect 134 -899 170 -843
rect -170 -1060 170 -899
rect -170 -1116 -134 -1060
rect -78 -1116 78 -1060
rect 134 -1116 170 -1060
rect -170 -1155 170 -1116
<< properties >>
string GDS_END 2266306
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2265022
<< end >>
