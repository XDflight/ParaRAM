magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -3793 23 3793 80
rect -3793 -23 -3739 23
rect -3693 -23 -3581 23
rect -3535 -23 -3423 23
rect -3377 -23 -3264 23
rect -3218 -23 -3106 23
rect -3060 -23 -2948 23
rect -2902 -23 -2790 23
rect -2744 -23 -2632 23
rect -2586 -23 -2474 23
rect -2428 -23 -2316 23
rect -2270 -23 -2158 23
rect -2112 -23 -2000 23
rect -1954 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1954 23
rect 2000 -23 2112 23
rect 2158 -23 2270 23
rect 2316 -23 2428 23
rect 2474 -23 2586 23
rect 2632 -23 2744 23
rect 2790 -23 2902 23
rect 2948 -23 3060 23
rect 3106 -23 3218 23
rect 3264 -23 3377 23
rect 3423 -23 3535 23
rect 3581 -23 3693 23
rect 3739 -23 3793 23
rect -3793 -80 3793 -23
<< psubdiffcont >>
rect -3739 -23 -3693 23
rect -3581 -23 -3535 23
rect -3423 -23 -3377 23
rect -3264 -23 -3218 23
rect -3106 -23 -3060 23
rect -2948 -23 -2902 23
rect -2790 -23 -2744 23
rect -2632 -23 -2586 23
rect -2474 -23 -2428 23
rect -2316 -23 -2270 23
rect -2158 -23 -2112 23
rect -2000 -23 -1954 23
rect -1841 -23 -1795 23
rect -1683 -23 -1637 23
rect -1525 -23 -1479 23
rect -1367 -23 -1321 23
rect -1209 -23 -1163 23
rect -1051 -23 -1005 23
rect -893 -23 -847 23
rect -735 -23 -689 23
rect -577 -23 -531 23
rect -418 -23 -372 23
rect -260 -23 -214 23
rect -102 -23 -56 23
rect 56 -23 102 23
rect 214 -23 260 23
rect 372 -23 418 23
rect 531 -23 577 23
rect 689 -23 735 23
rect 847 -23 893 23
rect 1005 -23 1051 23
rect 1163 -23 1209 23
rect 1321 -23 1367 23
rect 1479 -23 1525 23
rect 1637 -23 1683 23
rect 1795 -23 1841 23
rect 1954 -23 2000 23
rect 2112 -23 2158 23
rect 2270 -23 2316 23
rect 2428 -23 2474 23
rect 2586 -23 2632 23
rect 2744 -23 2790 23
rect 2902 -23 2948 23
rect 3060 -23 3106 23
rect 3218 -23 3264 23
rect 3377 -23 3423 23
rect 3535 -23 3581 23
rect 3693 -23 3739 23
<< metal1 >>
rect -3774 23 3774 60
rect -3774 -23 -3739 23
rect -3693 -23 -3581 23
rect -3535 -23 -3423 23
rect -3377 -23 -3264 23
rect -3218 -23 -3106 23
rect -3060 -23 -2948 23
rect -2902 -23 -2790 23
rect -2744 -23 -2632 23
rect -2586 -23 -2474 23
rect -2428 -23 -2316 23
rect -2270 -23 -2158 23
rect -2112 -23 -2000 23
rect -1954 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1954 23
rect 2000 -23 2112 23
rect 2158 -23 2270 23
rect 2316 -23 2428 23
rect 2474 -23 2586 23
rect 2632 -23 2744 23
rect 2790 -23 2902 23
rect 2948 -23 3060 23
rect 3106 -23 3218 23
rect 3264 -23 3377 23
rect 3423 -23 3535 23
rect 3581 -23 3693 23
rect 3739 -23 3774 23
rect -3774 -60 3774 -23
<< properties >>
string GDS_END 679126
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 675842
<< end >>
