magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< pwell >>
rect 5332 30656 28868 30688
rect 5332 -88 28868 -56
<< polysilicon >>
rect 5143 30529 5457 30548
rect 5143 30389 5162 30529
rect 5208 30394 5457 30529
rect 28741 30465 29111 30548
rect 28741 30419 28992 30465
rect 29038 30419 29111 30465
rect 28741 30394 29111 30419
rect 5208 30389 5227 30394
rect 5143 30370 5227 30389
rect 28919 30301 29111 30394
rect 28919 30255 28992 30301
rect 29038 30255 29111 30301
rect 28919 30209 29111 30255
rect 5143 28870 5457 29006
rect 5143 28730 5162 28870
rect 5208 28852 5457 28870
rect 28741 28905 29111 29006
rect 28741 28859 28992 28905
rect 29038 28859 29111 28905
rect 28741 28852 29111 28859
rect 5208 28748 5227 28852
rect 28919 28748 29111 28852
rect 5208 28730 5457 28748
rect 5143 28594 5457 28730
rect 28741 28741 29111 28748
rect 28741 28695 28992 28741
rect 29038 28695 29111 28741
rect 28741 28594 29111 28695
rect 5143 27070 5457 27206
rect 5143 26930 5162 27070
rect 5208 27052 5457 27070
rect 28741 27105 29111 27206
rect 28741 27059 28992 27105
rect 29038 27059 29111 27105
rect 28741 27052 29111 27059
rect 5208 26948 5227 27052
rect 28919 26948 29111 27052
rect 5208 26930 5457 26948
rect 5143 26794 5457 26930
rect 28741 26941 29111 26948
rect 28741 26895 28992 26941
rect 29038 26895 29111 26941
rect 28741 26794 29111 26895
rect 5143 25270 5457 25406
rect 5143 25130 5162 25270
rect 5208 25252 5457 25270
rect 28741 25305 29111 25406
rect 28741 25259 28992 25305
rect 29038 25259 29111 25305
rect 28741 25252 29111 25259
rect 5208 25148 5227 25252
rect 28919 25148 29111 25252
rect 5208 25130 5457 25148
rect 5143 24994 5457 25130
rect 28741 25141 29111 25148
rect 28741 25095 28992 25141
rect 29038 25095 29111 25141
rect 28741 24994 29111 25095
rect 5143 23470 5457 23606
rect 5143 23330 5162 23470
rect 5208 23452 5457 23470
rect 28741 23505 29111 23606
rect 28741 23459 28992 23505
rect 29038 23459 29111 23505
rect 28741 23452 29111 23459
rect 5208 23348 5227 23452
rect 28919 23348 29111 23452
rect 5208 23330 5457 23348
rect 5143 23194 5457 23330
rect 28741 23341 29111 23348
rect 28741 23295 28992 23341
rect 29038 23295 29111 23341
rect 28741 23194 29111 23295
rect 5143 21670 5457 21806
rect 5143 21530 5162 21670
rect 5208 21652 5457 21670
rect 28741 21705 29111 21806
rect 28741 21659 28992 21705
rect 29038 21659 29111 21705
rect 28741 21652 29111 21659
rect 5208 21548 5227 21652
rect 28919 21548 29111 21652
rect 5208 21530 5457 21548
rect 5143 21394 5457 21530
rect 28741 21541 29111 21548
rect 28741 21495 28992 21541
rect 29038 21495 29111 21541
rect 28741 21394 29111 21495
rect 5143 19870 5457 20006
rect 5143 19730 5162 19870
rect 5208 19852 5457 19870
rect 28741 19905 29111 20006
rect 28741 19859 28992 19905
rect 29038 19859 29111 19905
rect 28741 19852 29111 19859
rect 5208 19748 5227 19852
rect 28919 19748 29111 19852
rect 5208 19730 5457 19748
rect 5143 19594 5457 19730
rect 28741 19741 29111 19748
rect 28741 19695 28992 19741
rect 29038 19695 29111 19741
rect 28741 19594 29111 19695
rect 5143 18070 5457 18206
rect 5143 17930 5162 18070
rect 5208 18052 5457 18070
rect 28741 18105 29111 18206
rect 28741 18059 28992 18105
rect 29038 18059 29111 18105
rect 28741 18052 29111 18059
rect 5208 17948 5227 18052
rect 28919 17948 29111 18052
rect 5208 17930 5457 17948
rect 5143 17794 5457 17930
rect 28741 17941 29111 17948
rect 28741 17895 28992 17941
rect 29038 17895 29111 17941
rect 28741 17794 29111 17895
rect 5143 16270 5457 16406
rect 5143 16130 5162 16270
rect 5208 16252 5457 16270
rect 28741 16305 29111 16406
rect 28741 16259 28992 16305
rect 29038 16259 29111 16305
rect 28741 16252 29111 16259
rect 5208 16148 5227 16252
rect 28919 16148 29111 16252
rect 5208 16130 5457 16148
rect 5143 15994 5457 16130
rect 28741 16141 29111 16148
rect 28741 16095 28992 16141
rect 29038 16095 29111 16141
rect 28741 15994 29111 16095
rect 5143 14470 5457 14606
rect 5143 14330 5162 14470
rect 5208 14452 5457 14470
rect 28741 14505 29111 14606
rect 28741 14459 28992 14505
rect 29038 14459 29111 14505
rect 28741 14452 29111 14459
rect 5208 14348 5227 14452
rect 28919 14348 29111 14452
rect 5208 14330 5457 14348
rect 5143 14194 5457 14330
rect 28741 14341 29111 14348
rect 28741 14295 28992 14341
rect 29038 14295 29111 14341
rect 28741 14194 29111 14295
rect 5143 12670 5457 12806
rect 5143 12530 5162 12670
rect 5208 12652 5457 12670
rect 28741 12705 29111 12806
rect 28741 12659 28992 12705
rect 29038 12659 29111 12705
rect 28741 12652 29111 12659
rect 5208 12548 5227 12652
rect 28919 12548 29111 12652
rect 5208 12530 5457 12548
rect 5143 12394 5457 12530
rect 28741 12541 29111 12548
rect 28741 12495 28992 12541
rect 29038 12495 29111 12541
rect 28741 12394 29111 12495
rect 5143 10870 5457 11006
rect 5143 10730 5162 10870
rect 5208 10852 5457 10870
rect 28741 10905 29111 11006
rect 28741 10859 28992 10905
rect 29038 10859 29111 10905
rect 28741 10852 29111 10859
rect 5208 10748 5227 10852
rect 28919 10748 29111 10852
rect 5208 10730 5457 10748
rect 5143 10594 5457 10730
rect 28741 10741 29111 10748
rect 28741 10695 28992 10741
rect 29038 10695 29111 10741
rect 28741 10594 29111 10695
rect 5143 9070 5457 9206
rect 5143 8930 5162 9070
rect 5208 9052 5457 9070
rect 28741 9105 29111 9206
rect 28741 9059 28992 9105
rect 29038 9059 29111 9105
rect 28741 9052 29111 9059
rect 5208 8948 5227 9052
rect 28919 8948 29111 9052
rect 5208 8930 5457 8948
rect 5143 8794 5457 8930
rect 28741 8941 29111 8948
rect 28741 8895 28992 8941
rect 29038 8895 29111 8941
rect 28741 8794 29111 8895
rect 5143 7270 5457 7406
rect 5143 7130 5162 7270
rect 5208 7252 5457 7270
rect 28741 7305 29111 7406
rect 28741 7259 28992 7305
rect 29038 7259 29111 7305
rect 28741 7252 29111 7259
rect 5208 7148 5227 7252
rect 28919 7148 29111 7252
rect 5208 7130 5457 7148
rect 5143 6994 5457 7130
rect 28741 7141 29111 7148
rect 28741 7095 28992 7141
rect 29038 7095 29111 7141
rect 28741 6994 29111 7095
rect 5143 5470 5457 5606
rect 5143 5330 5162 5470
rect 5208 5452 5457 5470
rect 28741 5505 29111 5606
rect 28741 5459 28992 5505
rect 29038 5459 29111 5505
rect 28741 5452 29111 5459
rect 5208 5348 5227 5452
rect 28919 5348 29111 5452
rect 5208 5330 5457 5348
rect 5143 5194 5457 5330
rect 28741 5341 29111 5348
rect 28741 5295 28992 5341
rect 29038 5295 29111 5341
rect 28741 5194 29111 5295
rect 5143 3670 5457 3806
rect 5143 3530 5162 3670
rect 5208 3652 5457 3670
rect 28741 3705 29111 3806
rect 28741 3659 28992 3705
rect 29038 3659 29111 3705
rect 28741 3652 29111 3659
rect 5208 3548 5227 3652
rect 28919 3548 29111 3652
rect 5208 3530 5457 3548
rect 5143 3394 5457 3530
rect 28741 3541 29111 3548
rect 28741 3495 28992 3541
rect 29038 3495 29111 3541
rect 28741 3394 29111 3495
rect 5143 1870 5457 2006
rect 5143 1730 5162 1870
rect 5208 1852 5457 1870
rect 28741 1905 29111 2006
rect 28741 1859 28992 1905
rect 29038 1859 29111 1905
rect 28741 1852 29111 1859
rect 5208 1748 5227 1852
rect 28919 1748 29111 1852
rect 5208 1730 5457 1748
rect 5143 1594 5457 1730
rect 28741 1741 29111 1748
rect 28741 1695 28992 1741
rect 29038 1695 29111 1741
rect 28741 1594 29111 1695
rect 28919 345 29111 391
rect 28919 299 28992 345
rect 29038 299 29111 345
rect 5143 211 5227 230
rect 5143 71 5162 211
rect 5208 206 5227 211
rect 28919 206 29111 299
rect 5208 71 5457 206
rect 5143 52 5457 71
rect 28795 181 29111 206
rect 28795 135 28992 181
rect 29038 135 29111 181
rect 28795 52 29111 135
<< polycontact >>
rect 5162 30389 5208 30529
rect 28992 30419 29038 30465
rect 28992 30255 29038 30301
rect 5162 28730 5208 28870
rect 28992 28859 29038 28905
rect 28992 28695 29038 28741
rect 5162 26930 5208 27070
rect 28992 27059 29038 27105
rect 28992 26895 29038 26941
rect 5162 25130 5208 25270
rect 28992 25259 29038 25305
rect 28992 25095 29038 25141
rect 5162 23330 5208 23470
rect 28992 23459 29038 23505
rect 28992 23295 29038 23341
rect 5162 21530 5208 21670
rect 28992 21659 29038 21705
rect 28992 21495 29038 21541
rect 5162 19730 5208 19870
rect 28992 19859 29038 19905
rect 28992 19695 29038 19741
rect 5162 17930 5208 18070
rect 28992 18059 29038 18105
rect 28992 17895 29038 17941
rect 5162 16130 5208 16270
rect 28992 16259 29038 16305
rect 28992 16095 29038 16141
rect 5162 14330 5208 14470
rect 28992 14459 29038 14505
rect 28992 14295 29038 14341
rect 5162 12530 5208 12670
rect 28992 12659 29038 12705
rect 28992 12495 29038 12541
rect 5162 10730 5208 10870
rect 28992 10859 29038 10905
rect 28992 10695 29038 10741
rect 5162 8930 5208 9070
rect 28992 9059 29038 9105
rect 28992 8895 29038 8941
rect 5162 7130 5208 7270
rect 28992 7259 29038 7305
rect 28992 7095 29038 7141
rect 5162 5330 5208 5470
rect 28992 5459 29038 5505
rect 28992 5295 29038 5341
rect 5162 3530 5208 3670
rect 28992 3659 29038 3705
rect 28992 3495 29038 3541
rect 5162 1730 5208 1870
rect 28992 1859 29038 1905
rect 28992 1695 29038 1741
rect 28992 299 29038 345
rect 5162 71 5208 211
rect 28992 135 29038 181
<< metal1 >>
rect 5147 30529 5223 30540
rect 5147 30528 5162 30529
rect 5208 30528 5223 30529
rect 5147 30268 5159 30528
rect 5211 30268 5223 30528
rect 5147 30256 5223 30268
rect 28951 30470 29075 30510
rect 28951 30418 28987 30470
rect 29039 30418 29075 30470
rect 28951 30301 29075 30418
rect 28951 30255 28992 30301
rect 29038 30255 29075 30301
rect 28951 30252 29075 30255
rect 28951 30200 28987 30252
rect 29039 30200 29075 30252
rect 28951 30160 29075 30200
rect 5147 28930 5223 28942
rect 5147 28670 5159 28930
rect 5211 28670 5223 28930
rect 5147 28658 5223 28670
rect 28951 28933 29075 28973
rect 28951 28881 28987 28933
rect 29039 28881 29075 28933
rect 28951 28859 28992 28881
rect 29038 28859 29075 28881
rect 28951 28741 29075 28859
rect 28951 28715 28992 28741
rect 29038 28715 29075 28741
rect 28951 28663 28987 28715
rect 29039 28663 29075 28715
rect 28951 28623 29075 28663
rect 5147 27130 5223 27142
rect 5147 26870 5159 27130
rect 5211 26870 5223 27130
rect 5147 26858 5223 26870
rect 28951 27133 29075 27173
rect 28951 27081 28987 27133
rect 29039 27100 29075 27133
rect 29039 27081 29464 27100
rect 28951 27059 28992 27081
rect 29038 27059 29464 27081
rect 28951 26941 29464 27059
rect 28951 26915 28992 26941
rect 29038 26915 29464 26941
rect 28951 26863 28987 26915
rect 29039 26900 29464 26915
rect 29039 26863 29075 26900
rect 28951 26823 29075 26863
rect 5147 25330 5223 25342
rect 5147 25070 5159 25330
rect 5211 25070 5223 25330
rect 5147 25058 5223 25070
rect 28951 25337 29075 25377
rect 28951 25285 28987 25337
rect 29039 25285 29075 25337
rect 28951 25259 28992 25285
rect 29038 25259 29075 25285
rect 28951 25141 29075 25259
rect 28951 25119 28992 25141
rect 29038 25119 29075 25141
rect 28951 25067 28987 25119
rect 29039 25067 29075 25119
rect 28951 25027 29075 25067
rect 5143 23530 5219 23542
rect 5143 23270 5155 23530
rect 5207 23470 5219 23530
rect 5208 23330 5219 23470
rect 5207 23270 5219 23330
rect 5143 23258 5219 23270
rect 28951 23533 29075 23573
rect 28951 23481 28987 23533
rect 29039 23481 29075 23533
rect 28951 23459 28992 23481
rect 29038 23459 29075 23481
rect 28951 23341 29075 23459
rect 28951 23315 28992 23341
rect 29038 23315 29075 23341
rect 28951 23263 28987 23315
rect 29039 23263 29075 23315
rect 28951 23223 29075 23263
rect 5147 21730 5223 21742
rect 5147 21470 5159 21730
rect 5211 21470 5223 21730
rect 5147 21458 5223 21470
rect 28951 21737 29075 21777
rect 28951 21685 28987 21737
rect 29039 21685 29075 21737
rect 28951 21659 28992 21685
rect 29038 21659 29075 21685
rect 28951 21541 29075 21659
rect 28951 21519 28992 21541
rect 29038 21519 29075 21541
rect 28951 21467 28987 21519
rect 29039 21467 29075 21519
rect 28951 21427 29075 21467
rect 5147 19930 5223 19942
rect 5147 19670 5159 19930
rect 5211 19670 5223 19930
rect 5147 19658 5223 19670
rect 28951 19933 29075 19973
rect 28951 19881 28987 19933
rect 29039 19881 29075 19933
rect 28951 19859 28992 19881
rect 29038 19859 29075 19881
rect 28951 19741 29075 19859
rect 28951 19715 28992 19741
rect 29038 19715 29075 19741
rect 28951 19663 28987 19715
rect 29039 19663 29075 19715
rect 28951 19623 29075 19663
rect 5147 18130 5223 18142
rect 5147 17870 5159 18130
rect 5211 17870 5223 18130
rect 5147 17858 5223 17870
rect 28951 18137 29075 18177
rect 28951 18085 28987 18137
rect 29039 18085 29075 18137
rect 28951 18059 28992 18085
rect 29038 18059 29075 18085
rect 28951 17941 29075 18059
rect 28951 17919 28992 17941
rect 29038 17919 29075 17941
rect 28951 17867 28987 17919
rect 29039 17867 29075 17919
rect 28951 17827 29075 17867
rect 5147 16330 5223 16342
rect 5147 16070 5159 16330
rect 5211 16070 5223 16330
rect 5147 16058 5223 16070
rect 28951 16333 29075 16373
rect 28951 16281 28987 16333
rect 29039 16281 29075 16333
rect 28951 16259 28992 16281
rect 29038 16259 29075 16281
rect 28951 16141 29075 16259
rect 28951 16115 28992 16141
rect 29038 16115 29075 16141
rect 28951 16063 28987 16115
rect 29039 16063 29075 16115
rect 28951 16023 29075 16063
rect 5147 14530 5223 14542
rect 5147 14270 5159 14530
rect 5211 14270 5223 14530
rect 5147 14258 5223 14270
rect 28951 14537 29075 14577
rect 28951 14485 28987 14537
rect 29039 14485 29075 14537
rect 28951 14459 28992 14485
rect 29038 14459 29075 14485
rect 28951 14341 29075 14459
rect 28951 14319 28992 14341
rect 29038 14319 29075 14341
rect 28951 14267 28987 14319
rect 29039 14267 29075 14319
rect 28951 14227 29075 14267
rect 5147 12730 5223 12742
rect 5147 12470 5159 12730
rect 5211 12470 5223 12730
rect 5147 12458 5223 12470
rect 28951 12733 29075 12773
rect 28951 12681 28987 12733
rect 29039 12681 29075 12733
rect 28951 12659 28992 12681
rect 29038 12659 29075 12681
rect 28951 12541 29075 12659
rect 28951 12515 28992 12541
rect 29038 12515 29075 12541
rect 28951 12463 28987 12515
rect 29039 12463 29075 12515
rect 28951 12423 29075 12463
rect 5147 10930 5223 10942
rect 5147 10670 5159 10930
rect 5211 10670 5223 10930
rect 5147 10658 5223 10670
rect 28951 10937 29075 10977
rect 28951 10885 28987 10937
rect 29039 10885 29075 10937
rect 28951 10859 28992 10885
rect 29038 10859 29075 10885
rect 28951 10741 29075 10859
rect 28951 10719 28992 10741
rect 29038 10719 29075 10741
rect 28951 10667 28987 10719
rect 29039 10667 29075 10719
rect 28951 10627 29075 10667
rect 5147 9130 5223 9142
rect 5147 8870 5159 9130
rect 5211 8870 5223 9130
rect 5147 8858 5223 8870
rect 28951 9133 29075 9173
rect 28951 9081 28987 9133
rect 29039 9081 29075 9133
rect 28951 9059 28992 9081
rect 29038 9059 29075 9081
rect 28951 8941 29075 9059
rect 28951 8915 28992 8941
rect 29038 8915 29075 8941
rect 28951 8863 28987 8915
rect 29039 8863 29075 8915
rect 28951 8823 29075 8863
rect 5147 7330 5223 7342
rect 5147 7070 5159 7330
rect 5211 7070 5223 7330
rect 5147 7058 5223 7070
rect 28951 7337 29075 7377
rect 28951 7285 28987 7337
rect 29039 7285 29075 7337
rect 28951 7259 28992 7285
rect 29038 7259 29075 7285
rect 28951 7141 29075 7259
rect 28951 7119 28992 7141
rect 29038 7119 29075 7141
rect 28951 7067 28987 7119
rect 29039 7067 29075 7119
rect 28951 7027 29075 7067
rect 5147 5530 5223 5542
rect 5147 5270 5159 5530
rect 5211 5270 5223 5530
rect 5147 5258 5223 5270
rect 28951 5533 29075 5573
rect 28951 5481 28987 5533
rect 29039 5481 29075 5533
rect 28951 5459 28992 5481
rect 29038 5459 29075 5481
rect 28951 5341 29075 5459
rect 28951 5315 28992 5341
rect 29038 5315 29075 5341
rect 28951 5263 28987 5315
rect 29039 5263 29075 5315
rect 28951 5223 29075 5263
rect 5147 3730 5223 3742
rect 5147 3470 5159 3730
rect 5211 3470 5223 3730
rect 5147 3458 5223 3470
rect 28951 3737 29075 3777
rect 28951 3685 28987 3737
rect 29039 3685 29075 3737
rect 28951 3659 28992 3685
rect 29038 3659 29075 3685
rect 28951 3541 29075 3659
rect 28951 3519 28992 3541
rect 29038 3519 29075 3541
rect 28951 3467 28987 3519
rect 29039 3467 29075 3519
rect 28951 3427 29075 3467
rect 5147 1930 5223 1942
rect 5147 1670 5159 1930
rect 5211 1670 5223 1930
rect 5147 1658 5223 1670
rect 28951 1933 29075 1973
rect 28951 1881 28987 1933
rect 29039 1881 29075 1933
rect 28951 1859 28992 1881
rect 29038 1859 29075 1881
rect 28951 1741 29075 1859
rect 28951 1715 28992 1741
rect 29038 1715 29075 1741
rect 28951 1663 28987 1715
rect 29039 1663 29075 1715
rect 28951 1623 29075 1663
rect 28951 400 29075 440
rect 28951 348 28987 400
rect 29039 348 29075 400
rect 28951 345 29075 348
rect 28951 299 28992 345
rect 29038 299 29075 345
rect 5151 211 5219 222
rect 5151 71 5162 211
rect 5208 71 5219 211
rect 28951 182 29075 299
rect 28951 130 28987 182
rect 29039 130 29075 182
rect 28951 90 29075 130
rect 5151 60 5219 71
<< via1 >>
rect 5159 30389 5162 30528
rect 5162 30389 5208 30528
rect 5208 30389 5211 30528
rect 5159 30268 5211 30389
rect 28987 30465 29039 30470
rect 28987 30419 28992 30465
rect 28992 30419 29038 30465
rect 29038 30419 29039 30465
rect 28987 30418 29039 30419
rect 28987 30200 29039 30252
rect 5159 28870 5211 28930
rect 5159 28730 5162 28870
rect 5162 28730 5208 28870
rect 5208 28730 5211 28870
rect 5159 28670 5211 28730
rect 28987 28905 29039 28933
rect 28987 28881 28992 28905
rect 28992 28881 29038 28905
rect 29038 28881 29039 28905
rect 28987 28695 28992 28715
rect 28992 28695 29038 28715
rect 29038 28695 29039 28715
rect 28987 28663 29039 28695
rect 5159 27070 5211 27130
rect 5159 26930 5162 27070
rect 5162 26930 5208 27070
rect 5208 26930 5211 27070
rect 5159 26870 5211 26930
rect 28987 27105 29039 27133
rect 28987 27081 28992 27105
rect 28992 27081 29038 27105
rect 29038 27081 29039 27105
rect 28987 26895 28992 26915
rect 28992 26895 29038 26915
rect 29038 26895 29039 26915
rect 28987 26863 29039 26895
rect 5159 25270 5211 25330
rect 5159 25130 5162 25270
rect 5162 25130 5208 25270
rect 5208 25130 5211 25270
rect 5159 25070 5211 25130
rect 28987 25305 29039 25337
rect 28987 25285 28992 25305
rect 28992 25285 29038 25305
rect 29038 25285 29039 25305
rect 28987 25095 28992 25119
rect 28992 25095 29038 25119
rect 29038 25095 29039 25119
rect 28987 25067 29039 25095
rect 5155 23470 5207 23530
rect 5155 23330 5162 23470
rect 5162 23330 5207 23470
rect 5155 23270 5207 23330
rect 28987 23505 29039 23533
rect 28987 23481 28992 23505
rect 28992 23481 29038 23505
rect 29038 23481 29039 23505
rect 28987 23295 28992 23315
rect 28992 23295 29038 23315
rect 29038 23295 29039 23315
rect 28987 23263 29039 23295
rect 5159 21670 5211 21730
rect 5159 21530 5162 21670
rect 5162 21530 5208 21670
rect 5208 21530 5211 21670
rect 5159 21470 5211 21530
rect 28987 21705 29039 21737
rect 28987 21685 28992 21705
rect 28992 21685 29038 21705
rect 29038 21685 29039 21705
rect 28987 21495 28992 21519
rect 28992 21495 29038 21519
rect 29038 21495 29039 21519
rect 28987 21467 29039 21495
rect 5159 19870 5211 19930
rect 5159 19730 5162 19870
rect 5162 19730 5208 19870
rect 5208 19730 5211 19870
rect 5159 19670 5211 19730
rect 28987 19905 29039 19933
rect 28987 19881 28992 19905
rect 28992 19881 29038 19905
rect 29038 19881 29039 19905
rect 28987 19695 28992 19715
rect 28992 19695 29038 19715
rect 29038 19695 29039 19715
rect 28987 19663 29039 19695
rect 5159 18070 5211 18130
rect 5159 17930 5162 18070
rect 5162 17930 5208 18070
rect 5208 17930 5211 18070
rect 5159 17870 5211 17930
rect 28987 18105 29039 18137
rect 28987 18085 28992 18105
rect 28992 18085 29038 18105
rect 29038 18085 29039 18105
rect 28987 17895 28992 17919
rect 28992 17895 29038 17919
rect 29038 17895 29039 17919
rect 28987 17867 29039 17895
rect 5159 16270 5211 16330
rect 5159 16130 5162 16270
rect 5162 16130 5208 16270
rect 5208 16130 5211 16270
rect 5159 16070 5211 16130
rect 28987 16305 29039 16333
rect 28987 16281 28992 16305
rect 28992 16281 29038 16305
rect 29038 16281 29039 16305
rect 28987 16095 28992 16115
rect 28992 16095 29038 16115
rect 29038 16095 29039 16115
rect 28987 16063 29039 16095
rect 5159 14470 5211 14530
rect 5159 14330 5162 14470
rect 5162 14330 5208 14470
rect 5208 14330 5211 14470
rect 5159 14270 5211 14330
rect 28987 14505 29039 14537
rect 28987 14485 28992 14505
rect 28992 14485 29038 14505
rect 29038 14485 29039 14505
rect 28987 14295 28992 14319
rect 28992 14295 29038 14319
rect 29038 14295 29039 14319
rect 28987 14267 29039 14295
rect 5159 12670 5211 12730
rect 5159 12530 5162 12670
rect 5162 12530 5208 12670
rect 5208 12530 5211 12670
rect 5159 12470 5211 12530
rect 28987 12705 29039 12733
rect 28987 12681 28992 12705
rect 28992 12681 29038 12705
rect 29038 12681 29039 12705
rect 28987 12495 28992 12515
rect 28992 12495 29038 12515
rect 29038 12495 29039 12515
rect 28987 12463 29039 12495
rect 5159 10870 5211 10930
rect 5159 10730 5162 10870
rect 5162 10730 5208 10870
rect 5208 10730 5211 10870
rect 5159 10670 5211 10730
rect 28987 10905 29039 10937
rect 28987 10885 28992 10905
rect 28992 10885 29038 10905
rect 29038 10885 29039 10905
rect 28987 10695 28992 10719
rect 28992 10695 29038 10719
rect 29038 10695 29039 10719
rect 28987 10667 29039 10695
rect 5159 9070 5211 9130
rect 5159 8930 5162 9070
rect 5162 8930 5208 9070
rect 5208 8930 5211 9070
rect 5159 8870 5211 8930
rect 28987 9105 29039 9133
rect 28987 9081 28992 9105
rect 28992 9081 29038 9105
rect 29038 9081 29039 9105
rect 28987 8895 28992 8915
rect 28992 8895 29038 8915
rect 29038 8895 29039 8915
rect 28987 8863 29039 8895
rect 5159 7270 5211 7330
rect 5159 7130 5162 7270
rect 5162 7130 5208 7270
rect 5208 7130 5211 7270
rect 5159 7070 5211 7130
rect 28987 7305 29039 7337
rect 28987 7285 28992 7305
rect 28992 7285 29038 7305
rect 29038 7285 29039 7305
rect 28987 7095 28992 7119
rect 28992 7095 29038 7119
rect 29038 7095 29039 7119
rect 28987 7067 29039 7095
rect 5159 5470 5211 5530
rect 5159 5330 5162 5470
rect 5162 5330 5208 5470
rect 5208 5330 5211 5470
rect 5159 5270 5211 5330
rect 28987 5505 29039 5533
rect 28987 5481 28992 5505
rect 28992 5481 29038 5505
rect 29038 5481 29039 5505
rect 28987 5295 28992 5315
rect 28992 5295 29038 5315
rect 29038 5295 29039 5315
rect 28987 5263 29039 5295
rect 5159 3670 5211 3730
rect 5159 3530 5162 3670
rect 5162 3530 5208 3670
rect 5208 3530 5211 3670
rect 5159 3470 5211 3530
rect 28987 3705 29039 3737
rect 28987 3685 28992 3705
rect 28992 3685 29038 3705
rect 29038 3685 29039 3705
rect 28987 3495 28992 3519
rect 28992 3495 29038 3519
rect 29038 3495 29039 3519
rect 28987 3467 29039 3495
rect 5159 1870 5211 1930
rect 5159 1730 5162 1870
rect 5162 1730 5208 1870
rect 5208 1730 5211 1870
rect 5159 1670 5211 1730
rect 28987 1905 29039 1933
rect 28987 1881 28992 1905
rect 28992 1881 29038 1905
rect 29038 1881 29039 1905
rect 28987 1695 28992 1715
rect 28992 1695 29038 1715
rect 29038 1695 29039 1715
rect 28987 1663 29039 1695
rect 28987 348 29039 400
rect 28987 181 29039 182
rect 28987 135 28992 181
rect 28992 135 29038 181
rect 29038 135 29039 181
rect 28987 130 29039 135
<< metal2 >>
rect 5147 30528 5223 30540
rect 5147 30268 5159 30528
rect 5211 30268 5223 30528
rect 5147 28930 5223 30268
rect 5147 28670 5159 28930
rect 5211 28670 5223 28930
rect 5147 27130 5223 28670
rect 28950 30470 29075 30510
rect 28950 30418 28987 30470
rect 29039 30418 29075 30470
rect 28950 30252 29075 30418
rect 28950 30200 28987 30252
rect 29039 30200 29075 30252
rect 28950 28933 29075 30200
rect 28950 28881 28987 28933
rect 29039 28881 29075 28933
rect 28950 28715 29075 28881
rect 28950 28663 28987 28715
rect 29039 28663 29075 28715
rect 28950 28405 29075 28663
rect 5147 26870 5159 27130
rect 5211 26870 5223 27130
rect 5147 25330 5223 26870
rect 5147 25070 5159 25330
rect 5211 25070 5223 25330
rect 5147 23542 5223 25070
rect 5143 23530 5223 23542
rect 5143 23270 5155 23530
rect 5207 23270 5223 23530
rect 5143 23258 5223 23270
rect 5147 21730 5223 23258
rect 28950 27133 29075 27871
rect 28950 27081 28987 27133
rect 29039 27081 29075 27133
rect 28950 26915 29075 27081
rect 28950 26863 28987 26915
rect 29039 26863 29075 26915
rect 28950 25337 29075 26863
rect 28950 25285 28987 25337
rect 29039 25285 29075 25337
rect 28950 25119 29075 25285
rect 28950 25067 28987 25119
rect 29039 25067 29075 25119
rect 28950 23533 29075 25067
rect 28950 23481 28987 23533
rect 29039 23481 29075 23533
rect 28950 23315 29075 23481
rect 28950 23263 28987 23315
rect 29039 23263 29075 23315
rect 28950 22272 29075 23263
rect 5147 21470 5159 21730
rect 5211 21470 5223 21730
rect 5147 19930 5223 21470
rect 5147 19670 5159 19930
rect 5211 19670 5223 19930
rect 5147 18130 5223 19670
rect 5147 17870 5159 18130
rect 5211 17870 5223 18130
rect 5147 16330 5223 17870
rect 5147 16070 5159 16330
rect 5211 16070 5223 16330
rect 5147 14530 5223 16070
rect 5147 14270 5159 14530
rect 5211 14270 5223 14530
rect 5147 12730 5223 14270
rect 5147 12470 5159 12730
rect 5211 12470 5223 12730
rect 5147 10930 5223 12470
rect 5147 10670 5159 10930
rect 5211 10670 5223 10930
rect 5147 9130 5223 10670
rect 5147 8870 5159 9130
rect 5211 8870 5223 9130
rect 5147 7330 5223 8870
rect 5147 7070 5159 7330
rect 5211 7070 5223 7330
rect 5147 5530 5223 7070
rect 5147 5270 5159 5530
rect 5211 5270 5223 5530
rect 5147 3730 5223 5270
rect 5147 3470 5159 3730
rect 5211 3470 5223 3730
rect 5147 1930 5223 3470
rect 5147 1670 5159 1930
rect 5211 1670 5223 1930
rect 5147 134 5223 1670
rect 28950 21737 29075 21865
rect 28950 21685 28987 21737
rect 29039 21685 29075 21737
rect 28950 21519 29075 21685
rect 28950 21467 28987 21519
rect 29039 21467 29075 21519
rect 28950 19933 29075 21467
rect 28950 19881 28987 19933
rect 29039 19881 29075 19933
rect 28950 19715 29075 19881
rect 28950 19663 28987 19715
rect 29039 19663 29075 19715
rect 28950 18137 29075 19663
rect 28950 18085 28987 18137
rect 29039 18085 29075 18137
rect 28950 17919 29075 18085
rect 28950 17867 28987 17919
rect 29039 17867 29075 17919
rect 28950 16333 29075 17867
rect 28950 16281 28987 16333
rect 29039 16281 29075 16333
rect 28950 16115 29075 16281
rect 28950 16063 28987 16115
rect 29039 16063 29075 16115
rect 28950 14537 29075 16063
rect 28950 14485 28987 14537
rect 29039 14485 29075 14537
rect 28950 14319 29075 14485
rect 28950 14267 28987 14319
rect 29039 14267 29075 14319
rect 28950 12733 29075 14267
rect 28950 12681 28987 12733
rect 29039 12681 29075 12733
rect 28950 12515 29075 12681
rect 28950 12463 28987 12515
rect 29039 12463 29075 12515
rect 28950 10937 29075 12463
rect 28950 10885 28987 10937
rect 29039 10885 29075 10937
rect 28950 10719 29075 10885
rect 28950 10667 28987 10719
rect 29039 10667 29075 10719
rect 28950 9133 29075 10667
rect 28950 9081 28987 9133
rect 29039 9081 29075 9133
rect 28950 8915 29075 9081
rect 28950 8863 28987 8915
rect 29039 8863 29075 8915
rect 28950 7337 29075 8863
rect 28950 7285 28987 7337
rect 29039 7285 29075 7337
rect 28950 7119 29075 7285
rect 28950 7067 28987 7119
rect 29039 7067 29075 7119
rect 28950 5533 29075 7067
rect 28950 5481 28987 5533
rect 29039 5481 29075 5533
rect 28950 5315 29075 5481
rect 28950 5263 28987 5315
rect 29039 5263 29075 5315
rect 28950 3737 29075 5263
rect 28950 3685 28987 3737
rect 29039 3685 29075 3737
rect 28950 3519 29075 3685
rect 28950 3467 28987 3519
rect 29039 3467 29075 3519
rect 28950 1933 29075 3467
rect 28950 1881 28987 1933
rect 29039 1881 29075 1933
rect 28950 1715 29075 1881
rect 28950 1663 28987 1715
rect 29039 1663 29075 1715
rect 28950 400 29075 1663
rect 28950 348 28987 400
rect 29039 348 29075 400
rect 5147 -130 5157 134
rect 5213 -130 5223 134
rect 5147 -140 5223 -130
rect 28290 -786 28410 326
rect 28590 -786 28710 326
rect 28950 182 29075 348
rect 28950 130 28987 182
rect 29039 130 29075 182
rect 28950 90 29075 130
<< via2 >>
rect 5157 -130 5213 134
<< metal3 >>
rect 5147 134 5223 144
rect 5147 -130 5157 134
rect 5213 -130 5223 134
rect 5147 -140 5223 -130
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_0
timestamp 1666464484
transform -1 0 6000 0 1 20700
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_1
timestamp 1666464484
transform -1 0 6000 0 1 13500
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_2
timestamp 1666464484
transform -1 0 6000 0 1 2700
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_3
timestamp 1666464484
transform -1 0 6000 0 1 6300
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_4
timestamp 1666464484
transform -1 0 6000 0 1 18900
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_5
timestamp 1666464484
transform -1 0 6000 0 1 26100
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_6
timestamp 1666464484
transform -1 0 6000 0 1 11700
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_7
timestamp 1666464484
transform -1 0 6000 0 1 4500
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_8
timestamp 1666464484
transform -1 0 6000 0 1 8100
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_9
timestamp 1666464484
transform -1 0 6000 0 1 15300
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_10
timestamp 1666464484
transform -1 0 6000 0 1 22500
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_11
timestamp 1666464484
transform -1 0 6000 0 1 24300
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_12
timestamp 1666464484
transform -1 0 6000 0 1 17100
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_13
timestamp 1666464484
transform -1 0 6000 0 1 9900
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_14
timestamp 1666464484
transform -1 0 6000 0 1 27900
box -68 -68 668 1868
use 018SRAM_cell1_2x_256x8m81  018SRAM_cell1_2x_256x8m81_15
timestamp 1666464484
transform -1 0 6000 0 1 900
box -68 -68 668 1868
use 018SRAM_cell1_256x8m81  018SRAM_cell1_256x8m81_0
timestamp 1666464484
transform -1 0 6000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_256x8m81  018SRAM_cell1_256x8m81_1
timestamp 1666464484
transform -1 0 6000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_0
timestamp 1666464484
transform -1 0 22200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_1
timestamp 1666464484
transform -1 0 27000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_2
timestamp 1666464484
transform -1 0 26400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_3
timestamp 1666464484
transform -1 0 25800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_4
timestamp 1666464484
transform -1 0 25200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_5
timestamp 1666464484
transform -1 0 27600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_6
timestamp 1666464484
transform -1 0 24600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_7
timestamp 1666464484
transform -1 0 24000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_8
timestamp 1666464484
transform -1 0 23400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_9
timestamp 1666464484
transform -1 0 18000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_10
timestamp 1666464484
transform -1 0 18600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_11
timestamp 1666464484
transform -1 0 19800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_12
timestamp 1666464484
transform -1 0 19200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_13
timestamp 1666464484
transform -1 0 20400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_14
timestamp 1666464484
transform -1 0 21000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_15
timestamp 1666464484
transform -1 0 21600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_16
timestamp 1666464484
transform -1 0 8400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_17
timestamp 1666464484
transform -1 0 9600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_18
timestamp 1666464484
transform -1 0 10200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_19
timestamp 1666464484
transform -1 0 10800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_20
timestamp 1666464484
transform -1 0 11400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_21
timestamp 1666464484
transform -1 0 7200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_22
timestamp 1666464484
transform -1 0 16800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_23
timestamp 1666464484
transform -1 0 16200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_24
timestamp 1666464484
transform -1 0 15600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_25
timestamp 1666464484
transform -1 0 15000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_26
timestamp 1666464484
transform -1 0 13800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_27
timestamp 1666464484
transform -1 0 14400 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_28
timestamp 1666464484
transform -1 0 13200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_29
timestamp 1666464484
transform -1 0 12600 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_30
timestamp 1666464484
transform -1 0 7800 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_31
timestamp 1666464484
transform -1 0 9000 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_32
timestamp 1666464484
transform -1 0 12600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_33
timestamp 1666464484
transform -1 0 13200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_34
timestamp 1666464484
transform -1 0 14400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_35
timestamp 1666464484
transform -1 0 13800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_36
timestamp 1666464484
transform -1 0 15600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_37
timestamp 1666464484
transform -1 0 16200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_38
timestamp 1666464484
transform -1 0 16800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_39
timestamp 1666464484
transform -1 0 15000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_40
timestamp 1666464484
transform -1 0 7800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_41
timestamp 1666464484
transform -1 0 9000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_42
timestamp 1666464484
transform -1 0 8400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_43
timestamp 1666464484
transform -1 0 9600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_44
timestamp 1666464484
transform -1 0 10200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_45
timestamp 1666464484
transform -1 0 10800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_46
timestamp 1666464484
transform -1 0 11400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_47
timestamp 1666464484
transform -1 0 7200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_48
timestamp 1666464484
transform -1 0 18600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_49
timestamp 1666464484
transform -1 0 22200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_50
timestamp 1666464484
transform -1 0 21600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_51
timestamp 1666464484
transform -1 0 21000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_52
timestamp 1666464484
transform -1 0 20400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_53
timestamp 1666464484
transform -1 0 19200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_54
timestamp 1666464484
transform -1 0 19800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_55
timestamp 1666464484
transform -1 0 18000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_56
timestamp 1666464484
transform -1 0 27600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_57
timestamp 1666464484
transform -1 0 27000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_58
timestamp 1666464484
transform -1 0 26400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_59
timestamp 1666464484
transform -1 0 25800 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_60
timestamp 1666464484
transform -1 0 25200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_61
timestamp 1666464484
transform -1 0 24600 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_62
timestamp 1666464484
transform -1 0 24000 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_256x8m81  018SRAM_cell1_dummy_256x8m81_63
timestamp 1666464484
transform -1 0 23400 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_0
timestamp 1666464484
transform 1 0 28200 0 -1 1800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_1
timestamp 1666464484
transform 1 0 28200 0 1 0
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_2
timestamp 1666464484
transform 1 0 28200 0 -1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_3
timestamp 1666464484
transform 1 0 28200 0 -1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_4
timestamp 1666464484
transform 1 0 28200 0 -1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_5
timestamp 1666464484
transform 1 0 28200 0 -1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_6
timestamp 1666464484
transform 1 0 28200 0 -1 30600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_7
timestamp 1666464484
transform 1 0 28200 0 -1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_8
timestamp 1666464484
transform 1 0 28200 0 -1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_9
timestamp 1666464484
transform 1 0 28200 0 -1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_10
timestamp 1666464484
transform 1 0 28200 0 -1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_11
timestamp 1666464484
transform 1 0 28200 0 -1 18000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_12
timestamp 1666464484
transform 1 0 28200 0 -1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_13
timestamp 1666464484
transform 1 0 28200 0 -1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_14
timestamp 1666464484
transform 1 0 28200 0 -1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_15
timestamp 1666464484
transform 1 0 28200 0 -1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_16
timestamp 1666464484
transform 1 0 28200 0 -1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_17
timestamp 1666464484
transform 1 0 28200 0 -1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_18
timestamp 1666464484
transform 1 0 28200 0 1 5400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_19
timestamp 1666464484
transform 1 0 28200 0 1 7200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_20
timestamp 1666464484
transform 1 0 28200 0 1 10800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_21
timestamp 1666464484
transform 1 0 28200 0 1 14400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_22
timestamp 1666464484
transform 1 0 28200 0 1 18000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_23
timestamp 1666464484
transform 1 0 28200 0 1 21600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_24
timestamp 1666464484
transform 1 0 28200 0 1 25200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_25
timestamp 1666464484
transform 1 0 28200 0 1 28800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_26
timestamp 1666464484
transform 1 0 28200 0 1 3600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_27
timestamp 1666464484
transform 1 0 28200 0 1 9000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_28
timestamp 1666464484
transform 1 0 28200 0 1 12600
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_29
timestamp 1666464484
transform 1 0 28200 0 1 16200
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_30
timestamp 1666464484
transform 1 0 28200 0 1 19800
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_31
timestamp 1666464484
transform 1 0 28200 0 1 23400
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_32
timestamp 1666464484
transform 1 0 28200 0 1 27000
box -68 -68 668 968
use 018SRAM_cell1_dummy_R_256x8m81  018SRAM_cell1_dummy_R_256x8m81_33
timestamp 1666464484
transform 1 0 28200 0 1 1800
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_0
timestamp 1666464484
transform -1 0 22800 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_1
timestamp 1666464484
transform -1 0 12000 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_2
timestamp 1666464484
transform -1 0 6600 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_3
timestamp 1666464484
transform -1 0 12000 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_4
timestamp 1666464484
transform 1 0 27600 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_5
timestamp 1666464484
transform -1 0 22800 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_6
timestamp 1666464484
transform -1 0 17400 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_256x8m81  018SRAM_strap1_256x8m81_7
timestamp 1666464484
transform -1 0 17400 0 -1 30600
box -68 -68 668 968
use 018SRAM_strap1_bndry_256x8m81  018SRAM_strap1_bndry_256x8m81_0
timestamp 1666464484
transform 1 0 27600 0 1 0
box -68 -68 668 968
use 018SRAM_strap1_bndry_256x8m81  018SRAM_strap1_bndry_256x8m81_1
timestamp 1666464484
transform -1 0 6600 0 -1 30600
box -68 -68 668 968
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_0
timestamp 1666464484
transform 1 0 29015 0 -1 1800
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_1
timestamp 1666464484
transform 1 0 29015 0 -1 240
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_2
timestamp 1666464484
transform 1 0 29015 0 -1 3600
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_3
timestamp 1666464484
transform 1 0 29015 0 -1 27000
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_4
timestamp 1666464484
transform 1 0 29015 0 -1 23400
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_5
timestamp 1666464484
transform 1 0 29015 0 -1 19800
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_6
timestamp 1666464484
transform 1 0 29015 0 -1 28800
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_7
timestamp 1666464484
transform 1 0 29015 0 -1 25200
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_8
timestamp 1666464484
transform 1 0 29015 0 -1 21600
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_9
timestamp 1666464484
transform 1 0 29015 0 -1 16200
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_10
timestamp 1666464484
transform 1 0 29015 0 -1 12600
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_11
timestamp 1666464484
transform 1 0 29015 0 -1 9000
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_12
timestamp 1666464484
transform 1 0 29015 0 -1 18000
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_13
timestamp 1666464484
transform 1 0 29015 0 -1 14400
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_14
timestamp 1666464484
transform 1 0 29015 0 -1 10800
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_15
timestamp 1666464484
transform 1 0 29015 0 -1 7200
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_16
timestamp 1666464484
transform 1 0 29015 0 -1 5400
box 0 0 1 1
use M1_POLY2$$44754988_256x8m81  M1_POLY2$$44754988_256x8m81_17
timestamp 1666464484
transform 1 0 29015 0 -1 30360
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_0
timestamp 1666464484
transform 1 0 5185 0 1 1800
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_1
timestamp 1666464484
transform 1 0 5185 0 1 141
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_2
timestamp 1666464484
transform 1 0 5185 0 1 3600
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_3
timestamp 1666464484
transform 1 0 5185 0 1 7200
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_4
timestamp 1666464484
transform 1 0 5185 0 1 5400
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_5
timestamp 1666464484
transform 1 0 5185 0 1 14400
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_6
timestamp 1666464484
transform 1 0 5185 0 1 12600
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_7
timestamp 1666464484
transform 1 0 5185 0 1 16200
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_8
timestamp 1666464484
transform 1 0 5185 0 1 18000
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_9
timestamp 1666464484
transform 1 0 5185 0 1 21600
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_10
timestamp 1666464484
transform 1 0 5185 0 1 19800
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_11
timestamp 1666464484
transform 1 0 5185 0 1 23400
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_12
timestamp 1666464484
transform 1 0 5185 0 1 25200
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_13
timestamp 1666464484
transform 1 0 5185 0 1 28800
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_14
timestamp 1666464484
transform 1 0 5185 0 1 27000
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_15
timestamp 1666464484
transform 1 0 5185 0 1 30459
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_16
timestamp 1666464484
transform 1 0 5185 0 1 10800
box 0 0 1 1
use M1_POLY24310590878134_256x8m81  M1_POLY24310590878134_256x8m81_17
timestamp 1666464484
transform 1 0 5185 0 1 9000
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_0
timestamp 1666464484
transform 1 0 29013 0 -1 1798
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_1
timestamp 1666464484
transform 1 0 29013 0 -1 265
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_2
timestamp 1666464484
transform 1 0 29013 0 -1 23398
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_3
timestamp 1666464484
transform 1 0 29013 0 -1 19798
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_4
timestamp 1666464484
transform 1 0 29013 0 -1 16198
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_5
timestamp 1666464484
transform 1 0 29013 0 -1 12598
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_6
timestamp 1666464484
transform 1 0 29013 0 -1 8998
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_7
timestamp 1666464484
transform 1 0 29013 0 -1 5398
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_8
timestamp 1666464484
transform 1 0 29013 0 -1 10802
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_9
timestamp 1666464484
transform 1 0 29013 0 -1 25202
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_10
timestamp 1666464484
transform 1 0 29013 0 -1 18002
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_11
timestamp 1666464484
transform 1 0 29013 0 -1 3602
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_12
timestamp 1666464484
transform 1 0 29013 0 -1 14402
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_13
timestamp 1666464484
transform 1 0 29013 0 -1 28798
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_14
timestamp 1666464484
transform 1 0 29013 0 -1 21602
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_15
timestamp 1666464484
transform 1 0 29013 0 -1 7202
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_16
timestamp 1666464484
transform 1 0 29013 0 -1 30335
box 0 0 1 1
use M2_M1$$43375660_256x8m81  M2_M1$$43375660_256x8m81_17
timestamp 1666464484
transform 1 0 29013 0 -1 26998
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_0
timestamp 1666464484
transform 1 0 5185 0 1 1800
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_1
timestamp 1666464484
transform 1 0 5185 0 1 30398
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_2
timestamp 1666464484
transform 1 0 5185 0 1 28800
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_3
timestamp 1666464484
transform 1 0 5185 0 1 27000
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_4
timestamp 1666464484
transform 1 0 5185 0 1 25200
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_5
timestamp 1666464484
transform 1 0 5185 0 1 3600
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_6
timestamp 1666464484
transform 1 0 5185 0 1 5400
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_7
timestamp 1666464484
transform 1 0 5185 0 1 7200
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_8
timestamp 1666464484
transform 1 0 5185 0 1 9000
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_9
timestamp 1666464484
transform 1 0 5185 0 1 10800
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_10
timestamp 1666464484
transform 1 0 5185 0 1 12600
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_11
timestamp 1666464484
transform 1 0 5185 0 1 14400
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_12
timestamp 1666464484
transform 1 0 5185 0 1 16200
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_13
timestamp 1666464484
transform 1 0 5185 0 1 18000
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_14
timestamp 1666464484
transform 1 0 5185 0 1 19800
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_15
timestamp 1666464484
transform 1 0 5185 0 1 21600
box 0 0 1 1
use M2_M14310590878111_256x8m81  M2_M14310590878111_256x8m81_16
timestamp 1666464484
transform 1 0 5181 0 1 23400
box 0 0 1 1
use M3_M24310590878125_256x8m81  M3_M24310590878125_256x8m81_0
timestamp 1666464484
transform 1 0 5185 0 1 2
box 0 0 1 1
use rdummy_256x4_a_256x8m81  rdummy_256x4_a_256x8m81_0
timestamp 1666464484
transform 1 0 27562 0 1 -25410
box 0 0 1737 24714
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_0
timestamp 1666464484
transform -1 0 6600 0 1 27880
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_1
timestamp 1666464484
transform -1 0 6600 0 1 2680
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_2
timestamp 1666464484
transform -1 0 6600 0 1 4480
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_3
timestamp 1666464484
transform -1 0 6600 0 1 8080
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_4
timestamp 1666464484
transform -1 0 6600 0 1 6280
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_5
timestamp 1666464484
transform -1 0 6600 0 1 9880
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_6
timestamp 1666464484
transform -1 0 6600 0 1 11680
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_7
timestamp 1666464484
transform -1 0 6600 0 1 22480
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_8
timestamp 1666464484
transform -1 0 6600 0 1 24280
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_9
timestamp 1666464484
transform -1 0 6600 0 1 20680
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_10
timestamp 1666464484
transform -1 0 6600 0 1 18880
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_11
timestamp 1666464484
transform -1 0 6600 0 1 17080
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_12
timestamp 1666464484
transform -1 0 6600 0 1 15280
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_13
timestamp 1666464484
transform -1 0 6600 0 1 13480
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_14
timestamp 1666464484
transform -1 0 6600 0 1 26080
box -68 -48 668 1888
use strapx2b_bndry_256x8m81  strapx2b_bndry_256x8m81_15
timestamp 1666464484
transform -1 0 6600 0 1 880
box -68 -48 668 1888
<< labels >>
rlabel metal2 s 6302 880 6302 880 4 VDD
rlabel metal3 s 5934 29693 5934 29693 4 VDD
rlabel metal3 s 28266 1818 28266 1818 4 VSS
rlabel metal3 s 5934 1818 5934 1818 4 VSS
rlabel metal3 s 28266 893 28266 893 4 VDD
rlabel metal3 s 5934 893 5934 893 4 VDD
rlabel metal3 s 5562 30142 5562 30142 4 DWL
<< properties >>
string GDS_END 2068442
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2049752
<< end >>
