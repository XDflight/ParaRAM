magic
tech gf180mcuB
magscale 1 5
timestamp 1667403392
<< checkpaint >>
rect 6000 6000 36500 36500
<< metal4 >>
rect 7000 23034 8500 35500
tri 8500 23034 9122 23656 sw
tri 7000 21854 8180 23034 ne
rect 8180 21854 9122 23034
tri 9122 21854 10302 23034 sw
tri 8180 19732 10302 21854 ne
tri 10302 19732 12424 21854 sw
tri 10302 17610 12424 19732 ne
tri 12424 17610 14546 19732 sw
tri 12424 15488 14546 17610 ne
tri 14546 15488 16668 17610 sw
tri 14546 13366 16668 15488 ne
tri 16668 13366 18790 15488 sw
tri 16668 11244 18790 13366 ne
tri 18790 11244 20912 13366 sw
tri 18790 9122 20912 11244 ne
tri 20912 9122 23034 11244 sw
tri 20912 7000 23034 9122 ne
tri 23034 8500 23656 9122 sw
rect 23034 7000 35500 8500
<< end >>
