magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -802 28 803 66
rect -802 -28 -766 28
rect -710 -28 -555 28
rect -499 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 499 28
rect 555 -28 710 28
rect 766 -28 803 28
rect -802 -67 803 -28
<< via2 >>
rect -766 -28 -710 28
rect -555 -28 -499 28
rect -345 -28 -289 28
rect -134 -28 -78 28
rect 78 -28 134 28
rect 289 -28 345 28
rect 499 -28 555 28
rect 710 -28 766 28
<< metal3 >>
rect -803 28 803 67
rect -803 -28 -766 28
rect -710 -28 -555 28
rect -499 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 499 28
rect 555 -28 710 28
rect 766 -28 803 28
rect -803 -67 803 -28
<< properties >>
string GDS_END 577360
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 576716
<< end >>
