magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -19 354 19 360
rect -19 328 -13 354
rect 13 328 19 354
rect -19 292 19 328
rect -19 266 -13 292
rect 13 266 19 292
rect -19 230 19 266
rect -19 204 -13 230
rect 13 204 19 230
rect -19 168 19 204
rect -19 142 -13 168
rect 13 142 19 168
rect -19 106 19 142
rect -19 80 -13 106
rect 13 80 19 106
rect -19 44 19 80
rect -19 18 -13 44
rect 13 18 19 44
rect -19 -18 19 18
rect -19 -44 -13 -18
rect 13 -44 19 -18
rect -19 -80 19 -44
rect -19 -106 -13 -80
rect 13 -106 19 -80
rect -19 -142 19 -106
rect -19 -168 -13 -142
rect 13 -168 19 -142
rect -19 -204 19 -168
rect -19 -230 -13 -204
rect 13 -230 19 -204
rect -19 -266 19 -230
rect -19 -292 -13 -266
rect 13 -292 19 -266
rect -19 -328 19 -292
rect -19 -354 -13 -328
rect 13 -354 19 -328
rect -19 -360 19 -354
<< via1 >>
rect -13 328 13 354
rect -13 266 13 292
rect -13 204 13 230
rect -13 142 13 168
rect -13 80 13 106
rect -13 18 13 44
rect -13 -44 13 -18
rect -13 -106 13 -80
rect -13 -168 13 -142
rect -13 -230 13 -204
rect -13 -292 13 -266
rect -13 -354 13 -328
<< metal2 >>
rect -19 354 19 360
rect -19 328 -13 354
rect 13 328 19 354
rect -19 292 19 328
rect -19 266 -13 292
rect 13 266 19 292
rect -19 230 19 266
rect -19 204 -13 230
rect 13 204 19 230
rect -19 168 19 204
rect -19 142 -13 168
rect 13 142 19 168
rect -19 106 19 142
rect -19 80 -13 106
rect 13 80 19 106
rect -19 44 19 80
rect -19 18 -13 44
rect 13 18 19 44
rect -19 -18 19 18
rect -19 -44 -13 -18
rect 13 -44 19 -18
rect -19 -80 19 -44
rect -19 -106 -13 -80
rect 13 -106 19 -80
rect -19 -142 19 -106
rect -19 -168 -13 -142
rect 13 -168 19 -142
rect -19 -204 19 -168
rect -19 -230 -13 -204
rect 13 -230 19 -204
rect -19 -266 19 -230
rect -19 -292 -13 -266
rect 13 -292 19 -266
rect -19 -328 19 -292
rect -19 -354 -13 -328
rect 13 -354 19 -328
rect -19 -360 19 -354
<< properties >>
string GDS_END 634088
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 633188
<< end >>
