magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 766
<< polysilicon >>
rect -31 3538 88 3610
rect -31 -73 88 0
use pmos_5p04310590548768_128x8m81  pmos_5p04310590548768_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 3658
<< properties >>
string GDS_END 274654
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 274340
<< end >>
