magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 6048 844
rect 326 626 372 724
rect 1280 689 1348 724
rect 1963 620 2009 724
rect 74 354 318 430
rect 923 354 1695 430
rect 2404 518 2472 724
rect 2812 518 2880 724
rect 3234 518 3302 724
rect 3489 572 3535 676
rect 3693 646 3739 724
rect 3917 572 3963 676
rect 4141 646 4187 724
rect 4365 572 4411 676
rect 4589 646 4635 724
rect 4793 572 4839 676
rect 4997 646 5043 724
rect 5201 572 5247 676
rect 5405 646 5451 724
rect 5609 572 5656 676
rect 3489 492 5656 572
rect 5813 506 5859 724
rect 4608 253 4688 492
rect 283 60 329 152
rect 1230 60 1302 95
rect 1854 60 1926 95
rect 2359 60 2405 186
rect 2807 60 2853 186
rect 4150 227 5322 253
rect 3255 60 3301 186
rect 3424 173 5776 227
rect 3692 60 3760 127
rect 4140 60 4208 127
rect 4588 60 4656 127
rect 5036 60 5104 127
rect 5445 60 5552 127
rect 5943 60 5989 183
rect 0 -60 6048 60
<< obsm1 >>
rect 122 573 168 676
rect 519 643 1234 671
rect 1394 643 1898 671
rect 519 625 1898 643
rect 826 602 1898 625
rect 122 514 433 573
rect 387 464 433 514
rect 387 418 675 464
rect 387 245 433 418
rect 734 372 780 578
rect 59 198 433 245
rect 605 326 780 372
rect 59 143 105 198
rect 605 177 651 326
rect 826 280 872 602
rect 1188 597 1440 602
rect 1852 568 1898 602
rect 2211 568 2257 676
rect 1030 551 1133 556
rect 1486 551 1800 556
rect 1030 505 1800 551
rect 1852 522 2257 568
rect 1754 380 1800 505
rect 2211 472 2257 522
rect 2619 472 2665 676
rect 3027 472 3073 676
rect 2211 439 3301 472
rect 2211 426 4530 439
rect 3255 392 4530 426
rect 762 198 872 280
rect 1754 330 3193 380
rect 1754 279 1800 330
rect 3255 284 4095 319
rect 918 233 1800 279
rect 2211 273 4095 284
rect 2211 238 3301 273
rect 4881 392 5768 439
rect 5372 273 5897 319
rect 918 198 990 233
rect 1542 198 1614 233
rect 2211 187 2257 238
rect 507 152 651 177
rect 1138 152 1431 187
rect 1711 152 2257 187
rect 507 141 2257 152
rect 507 106 1184 141
rect 1385 106 1757 141
rect 2583 116 2629 238
rect 3031 116 3077 238
<< labels >>
rlabel metal1 s 74 354 318 430 6 EN
port 1 nsew default input
rlabel metal1 s 923 354 1695 430 6 I
port 2 nsew default input
rlabel metal1 s 5609 572 5656 676 6 ZN
port 3 nsew default output
rlabel metal1 s 5201 572 5247 676 6 ZN
port 3 nsew default output
rlabel metal1 s 4793 572 4839 676 6 ZN
port 3 nsew default output
rlabel metal1 s 4365 572 4411 676 6 ZN
port 3 nsew default output
rlabel metal1 s 3917 572 3963 676 6 ZN
port 3 nsew default output
rlabel metal1 s 3489 572 3535 676 6 ZN
port 3 nsew default output
rlabel metal1 s 3489 492 5656 572 6 ZN
port 3 nsew default output
rlabel metal1 s 4608 253 4688 492 6 ZN
port 3 nsew default output
rlabel metal1 s 4150 227 5322 253 6 ZN
port 3 nsew default output
rlabel metal1 s 3424 173 5776 227 6 ZN
port 3 nsew default output
rlabel metal1 s 0 724 6048 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 689 5859 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5405 689 5451 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4997 689 5043 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4589 689 4635 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4141 689 4187 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3693 689 3739 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 689 3302 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 689 2880 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 689 2472 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 689 2009 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1280 689 1348 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 689 372 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 646 5859 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5405 646 5451 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4997 646 5043 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4589 646 4635 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4141 646 4187 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3693 646 3739 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 646 3302 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 646 2880 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 646 2472 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 646 2009 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 646 372 689 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 626 5859 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 626 3302 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 626 2880 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 626 2472 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 626 2009 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 626 372 646 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 620 5859 626 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 620 3302 626 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 620 2880 626 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 620 2472 626 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1963 620 2009 626 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 518 5859 620 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3234 518 3302 620 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2812 518 2880 620 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2404 518 2472 620 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5813 506 5859 518 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3255 183 3301 186 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2807 183 2853 186 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2359 183 2405 186 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5943 152 5989 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3255 152 3301 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2807 152 2853 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2359 152 2405 183 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5943 127 5989 152 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3255 127 3301 152 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2807 127 2853 152 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2359 127 2405 152 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 283 127 329 152 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5943 95 5989 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5445 95 5552 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5036 95 5104 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4588 95 4656 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 95 4208 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3692 95 3760 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3255 95 3301 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2807 95 2853 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2359 95 2405 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 283 95 329 127 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5943 60 5989 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5445 60 5552 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5036 60 5104 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4588 60 4656 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 60 4208 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3692 60 3760 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3255 60 3301 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2807 60 2853 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2359 60 2405 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1854 60 1926 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1230 60 1302 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 283 60 329 95 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 6048 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 6048 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 553708
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 540842
<< end >>
