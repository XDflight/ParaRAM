magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 534 870
<< pwell >>
rect -86 -86 534 352
<< mvnmos >>
rect 125 68 245 232
<< mvpmos >>
rect 125 472 225 716
<< mvndiff >>
rect 37 172 125 232
rect 37 126 50 172
rect 96 126 125 172
rect 37 68 125 126
rect 245 175 333 232
rect 245 129 274 175
rect 320 129 333 175
rect 245 68 333 129
<< mvpdiff >>
rect 37 649 125 716
rect 37 509 50 649
rect 96 509 125 649
rect 37 472 125 509
rect 225 649 313 716
rect 225 509 254 649
rect 300 509 313 649
rect 225 472 313 509
<< mvndiffc >>
rect 50 126 96 172
rect 274 129 320 175
<< mvpdiffc >>
rect 50 509 96 649
rect 254 509 300 649
<< polysilicon >>
rect 125 716 225 760
rect 125 327 225 472
rect 125 314 245 327
rect 125 268 186 314
rect 232 268 245 314
rect 125 232 245 268
rect 125 24 245 68
<< polycontact >>
rect 186 268 232 314
<< metal1 >>
rect 0 724 448 844
rect 50 649 96 724
rect 50 472 96 509
rect 244 649 316 678
rect 244 509 254 649
rect 300 509 316 649
rect 244 461 316 509
rect 175 268 186 314
rect 232 268 320 314
rect 175 267 320 268
rect 50 172 96 232
rect 50 60 96 126
rect 274 175 320 267
rect 274 106 320 129
rect 0 -60 448 60
<< labels >>
flabel metal1 s 244 461 316 678 0 FreeSans 400 0 0 0 Z
port 1 nsew default output
flabel metal1 s 0 724 448 844 0 FreeSans 400 0 0 0 VDD
port 2 nsew power bidirectional abutment
flabel metal1 s 50 60 96 232 0 FreeSans 400 0 0 0 VSS
port 5 nsew ground bidirectional abutment
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 50 472 96 724 1 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 -60 448 60 1 VSS
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string GDS_END 312146
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 310188
string LEFclass core TIEHIGH
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
