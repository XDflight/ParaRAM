magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 254 -148 3069 1110
rect 4720 -71 7235 1078
rect 8460 -92 9060 1128
rect 14258 901 18305 1127
rect 23621 1109 24063 1110
rect 14258 -1 19596 901
rect 14258 -71 18226 -1
rect 21248 -4 24063 1109
rect 23621 -148 24063 -4
<< nmos >>
rect 13291 717 13921 837
rect 3267 248 4267 368
rect 13291 504 13921 624
rect 13291 280 13921 400
rect 20050 248 21050 368
<< ndiff >>
rect 13291 923 13921 969
rect 13291 877 13335 923
rect 13381 877 13502 923
rect 13548 877 13667 923
rect 13713 877 13832 923
rect 13878 877 13921 923
rect 13291 837 13921 877
rect 13291 624 13921 717
rect 3267 368 4267 493
rect 3267 216 4267 248
rect 3267 170 3412 216
rect 3458 170 3598 216
rect 3644 170 3785 216
rect 3831 170 3972 216
rect 4018 170 4158 216
rect 4204 170 4267 216
rect 13291 400 13921 504
rect 13291 230 13921 280
rect 3267 124 4267 170
rect 13291 184 13335 230
rect 13381 184 13502 230
rect 13548 184 13667 230
rect 13713 184 13832 230
rect 13878 184 13921 230
rect 20050 368 21050 493
rect 20050 216 21050 248
rect 13291 137 13921 184
rect 20050 170 20112 216
rect 20158 170 20299 216
rect 20345 170 20486 216
rect 20532 170 20672 216
rect 20718 170 20859 216
rect 20905 170 21050 216
rect 20050 124 21050 170
<< ndiffc >>
rect 13335 877 13381 923
rect 13502 877 13548 923
rect 13667 877 13713 923
rect 13832 877 13878 923
rect 3412 170 3458 216
rect 3598 170 3644 216
rect 3785 170 3831 216
rect 3972 170 4018 216
rect 4158 170 4204 216
rect 13335 184 13381 230
rect 13502 184 13548 230
rect 13667 184 13713 230
rect 13832 184 13878 230
rect 20112 170 20158 216
rect 20299 170 20345 216
rect 20486 170 20532 216
rect 20672 170 20718 216
rect 20859 170 20905 216
<< psubdiff >>
rect 7534 923 8088 942
rect 7534 877 7553 923
rect 8069 877 8088 923
rect 7534 858 8088 877
rect 4457 23 4613 80
rect 4457 -23 4512 23
rect 4558 -23 4613 23
rect 4457 -80 4613 -23
rect 19699 23 19859 83
rect 19699 -23 19756 23
rect 19802 -23 19859 23
rect 19699 -83 19859 -23
<< nsubdiff >>
rect 396 799 552 962
rect 5944 923 6457 969
rect 5944 877 6085 923
rect 6319 877 6457 923
rect 396 753 451 799
rect 497 753 552 799
rect 396 635 552 753
rect 5944 831 6457 877
rect 8603 923 8917 980
rect 15160 969 18162 980
rect 8603 877 8658 923
rect 8704 877 8816 923
rect 8862 877 8917 923
rect 8603 820 8917 877
rect 396 589 451 635
rect 497 589 552 635
rect 396 472 552 589
rect 396 426 451 472
rect 497 426 552 472
rect 396 309 552 426
rect 396 263 451 309
rect 497 263 552 309
rect 15160 923 18305 969
rect 15160 877 15215 923
rect 15261 877 15373 923
rect 15419 877 15531 923
rect 15577 877 15689 923
rect 15735 877 15847 923
rect 15893 877 16005 923
rect 16051 877 16164 923
rect 16210 877 16322 923
rect 16368 877 16480 923
rect 16526 877 16638 923
rect 16684 877 16796 923
rect 16842 877 16954 923
rect 17000 877 17112 923
rect 17158 877 17271 923
rect 17317 877 17429 923
rect 17475 877 17587 923
rect 17633 877 17745 923
rect 17791 877 17903 923
rect 17949 877 18061 923
rect 18107 901 18305 923
rect 18107 877 18362 901
rect 15160 831 18362 877
rect 15160 759 18162 831
rect 15160 713 15215 759
rect 15261 713 15373 759
rect 15419 713 15531 759
rect 15577 713 15689 759
rect 15735 713 15847 759
rect 15893 713 16005 759
rect 16051 713 16164 759
rect 16210 713 16322 759
rect 16368 713 16480 759
rect 16526 713 16638 759
rect 16684 713 16796 759
rect 16842 713 16954 759
rect 17000 713 17112 759
rect 17158 713 17271 759
rect 17317 713 17429 759
rect 17475 713 17587 759
rect 17633 713 17745 759
rect 17791 713 17903 759
rect 17949 713 18061 759
rect 18107 713 18162 759
rect 23764 799 23920 962
rect 23764 753 23819 799
rect 23865 753 23920 799
rect 15160 656 18162 713
rect 396 146 552 263
rect 396 100 451 146
rect 497 100 552 146
rect 23764 635 23920 753
rect 23764 589 23819 635
rect 23865 589 23920 635
rect 23764 146 23920 589
rect 396 -1 552 100
rect 23764 100 23819 146
rect 23865 100 23920 146
rect 23764 -1 23920 100
<< psubdiffcont >>
rect 7553 877 8069 923
rect 4512 -23 4558 23
rect 19756 -23 19802 23
<< nsubdiffcont >>
rect 6085 877 6319 923
rect 451 753 497 799
rect 8658 877 8704 923
rect 8816 877 8862 923
rect 451 589 497 635
rect 451 426 497 472
rect 451 263 497 309
rect 15215 877 15261 923
rect 15373 877 15419 923
rect 15531 877 15577 923
rect 15689 877 15735 923
rect 15847 877 15893 923
rect 16005 877 16051 923
rect 16164 877 16210 923
rect 16322 877 16368 923
rect 16480 877 16526 923
rect 16638 877 16684 923
rect 16796 877 16842 923
rect 16954 877 17000 923
rect 17112 877 17158 923
rect 17271 877 17317 923
rect 17429 877 17475 923
rect 17587 877 17633 923
rect 17745 877 17791 923
rect 17903 877 17949 923
rect 18061 877 18107 923
rect 15215 713 15261 759
rect 15373 713 15419 759
rect 15531 713 15577 759
rect 15689 713 15735 759
rect 15847 713 15893 759
rect 16005 713 16051 759
rect 16164 713 16210 759
rect 16322 713 16368 759
rect 16480 713 16526 759
rect 16638 713 16684 759
rect 16796 713 16842 759
rect 16954 713 17000 759
rect 17112 713 17158 759
rect 17271 713 17317 759
rect 17429 713 17475 759
rect 17587 713 17633 759
rect 17745 713 17791 759
rect 17903 713 17949 759
rect 18061 713 18107 759
rect 23819 753 23865 799
rect 451 100 497 146
rect 23819 589 23865 635
rect 23819 100 23865 146
<< polysilicon >>
rect 2968 757 3368 848
rect 2968 728 3091 757
rect 3072 624 3091 728
rect 2961 504 3091 624
rect 3054 400 3091 504
rect 2961 335 3091 400
rect 3137 728 3368 757
rect 9758 728 9942 848
rect 14047 837 14989 848
rect 3137 624 3156 728
rect 9858 710 9942 728
rect 12950 782 13291 837
rect 12950 736 12969 782
rect 13109 736 13291 782
rect 12950 717 13291 736
rect 13921 728 14989 837
rect 13921 717 14148 728
rect 9858 664 9877 710
rect 9923 664 9942 710
rect 9858 645 9942 664
rect 21047 728 21384 848
rect 21152 727 21261 728
rect 21152 624 21196 727
rect 3137 504 3368 624
rect 3137 335 3156 504
rect 4729 368 4788 537
rect 2961 280 3156 335
rect 3216 248 3267 368
rect 4267 248 4788 368
rect 4729 193 4788 248
rect 6027 438 6136 537
rect 6027 298 6071 438
rect 6117 298 6136 438
rect 6027 193 6136 298
rect 6274 438 6369 537
rect 6274 298 6293 438
rect 6339 298 6369 438
rect 7422 417 7492 537
rect 8153 440 8330 537
rect 13221 504 13291 624
rect 13921 587 14394 624
rect 13921 541 13954 587
rect 14094 541 14394 587
rect 13921 504 14394 541
rect 8153 417 8265 440
rect 8223 313 8265 417
rect 6274 193 6369 298
rect 7422 193 7492 313
rect 8153 300 8265 313
rect 8311 300 8330 440
rect 18199 465 18301 537
rect 8153 193 8330 300
rect 8535 279 9505 313
rect 13221 280 13291 400
rect 13921 356 15219 400
rect 13921 310 15060 356
rect 15200 310 15219 356
rect 13921 280 15219 310
rect 18199 325 18218 465
rect 18264 325 18301 465
rect 8535 233 9440 279
rect 9486 233 9505 279
rect 8535 193 9505 233
rect 18199 193 18301 325
rect 19528 368 19587 537
rect 21079 504 21196 624
rect 19528 248 20050 368
rect 21050 248 21094 368
rect 21177 305 21196 504
rect 21242 624 21261 727
rect 21242 504 21384 624
rect 21242 400 21263 504
rect 21242 305 21384 400
rect 21177 280 21384 305
rect 19528 193 19587 248
<< polycontact >>
rect 3091 335 3137 757
rect 12969 736 13109 782
rect 9877 664 9923 710
rect 6071 298 6117 438
rect 6293 298 6339 438
rect 13954 541 14094 587
rect 8265 300 8311 440
rect 15060 310 15200 356
rect 18218 325 18264 465
rect 9440 233 9486 279
rect 21196 305 21242 727
<< metal1 >>
rect 344 799 636 967
rect 3843 960 4604 966
rect 3842 926 4604 960
rect 3842 874 3880 926
rect 3932 874 4091 926
rect 4143 874 4303 926
rect 4355 874 4514 926
rect 4566 874 4604 926
rect 3842 840 4604 874
rect 3843 833 4604 840
rect 4778 960 5960 967
rect 7542 966 7920 967
rect 4778 926 6554 960
rect 4778 874 4816 926
rect 4868 874 5026 926
rect 5078 874 5237 926
rect 5289 874 5449 926
rect 5501 874 5660 926
rect 5712 874 5870 926
rect 5922 923 6554 926
rect 5922 877 6085 923
rect 6319 877 6554 923
rect 5922 874 6554 877
rect 4778 840 6554 874
rect 7542 926 8438 966
rect 7542 923 7926 926
rect 7978 923 8137 926
rect 7542 877 7553 923
rect 8069 877 8137 923
rect 7542 874 7926 877
rect 7978 874 8137 877
rect 8189 874 8348 926
rect 8400 874 8438 926
rect 4778 833 5960 840
rect 7542 833 8438 874
rect 8610 960 8918 967
rect 9811 960 10119 967
rect 13349 960 14110 966
rect 8610 926 8919 960
rect 8610 874 8648 926
rect 8700 923 8828 926
rect 8704 877 8816 923
rect 8700 874 8828 877
rect 8880 874 8919 926
rect 344 753 451 799
rect 497 753 636 799
rect 344 635 636 753
rect 3080 757 3148 768
rect 344 589 451 635
rect 497 589 636 635
rect 2615 702 2923 743
rect 2615 650 2653 702
rect 2705 650 2833 702
rect 2885 650 2923 702
rect 2615 610 2923 650
rect 344 497 636 589
rect 344 472 1089 497
rect 344 426 451 472
rect 497 426 1089 472
rect 344 378 1089 426
rect 344 309 636 378
rect 344 263 451 309
rect 497 263 636 309
rect 3080 335 3091 757
rect 3137 335 3148 757
rect 3377 710 3685 751
rect 3377 658 3415 710
rect 3467 658 3595 710
rect 3647 658 3685 710
rect 3377 618 3685 658
rect 4890 624 5862 664
rect 7449 661 7757 677
rect 4890 572 4928 624
rect 4980 572 5139 624
rect 5191 572 5350 624
rect 5402 572 5561 624
rect 5613 572 5772 624
rect 5824 572 5862 624
rect 4890 532 5862 572
rect 6034 541 6549 661
rect 7035 636 7757 661
rect 7035 584 7487 636
rect 7539 584 7667 636
rect 7719 584 7757 636
rect 7035 544 7757 584
rect 7035 541 7527 544
rect 3824 464 4314 504
rect 3824 412 3863 464
rect 3915 412 4043 464
rect 4095 412 4223 464
rect 4275 412 4314 464
rect 6034 438 6150 541
rect 3824 371 4314 412
rect 344 146 636 263
rect 2615 254 2923 295
rect 2615 202 2653 254
rect 2705 202 2833 254
rect 2885 202 2923 254
rect 2615 162 2923 202
rect 3080 253 3148 335
rect 4560 310 5956 432
rect 4560 253 4678 310
rect 3080 216 4678 253
rect 3080 170 3412 216
rect 3458 170 3598 216
rect 3644 170 3785 216
rect 3831 170 3972 216
rect 4018 170 4158 216
rect 4204 170 4678 216
rect 6034 298 6071 438
rect 6117 298 6150 438
rect 3080 162 4678 170
rect 4890 164 5862 204
rect 344 100 451 146
rect 497 100 636 146
rect 3080 133 4239 162
rect 344 -67 636 100
rect 4890 112 4928 164
rect 4980 112 5139 164
rect 5191 112 5350 164
rect 5402 112 5561 164
rect 5613 112 5772 164
rect 5824 112 5862 164
rect 4466 67 4621 74
rect 4890 72 5862 112
rect 6034 198 6150 298
rect 6236 438 6369 461
rect 6236 389 6293 438
rect 6236 337 6274 389
rect 6236 298 6293 337
rect 6339 298 6369 438
rect 8254 440 8322 451
rect 6520 430 7281 436
rect 6519 429 7281 430
rect 6519 396 7527 429
rect 6519 344 6557 396
rect 6609 344 6768 396
rect 6820 344 6980 396
rect 7032 344 7191 396
rect 7243 344 7527 396
rect 6519 310 7527 344
rect 6520 303 7281 310
rect 6236 278 6369 298
rect 8254 300 8265 440
rect 8311 300 8322 440
rect 8610 310 8919 874
rect 9088 926 10698 960
rect 13300 937 14110 960
rect 9088 874 9849 926
rect 9901 874 10029 926
rect 10081 874 10698 926
rect 9088 840 10698 874
rect 11888 926 14110 937
rect 11888 923 13386 926
rect 11888 877 13335 923
rect 13381 877 13386 923
rect 11888 874 13386 877
rect 13438 923 13597 926
rect 13438 877 13502 923
rect 13548 877 13597 923
rect 13438 874 13597 877
rect 13649 923 13809 926
rect 13861 923 14020 926
rect 13649 877 13667 923
rect 13713 877 13809 923
rect 13878 877 14020 923
rect 13649 874 13809 877
rect 13861 874 14020 877
rect 14072 874 14110 926
rect 11888 863 14110 874
rect 13300 840 14110 863
rect 9088 310 9204 840
rect 9811 834 10119 840
rect 13349 833 14110 840
rect 14392 960 14942 966
rect 18396 960 19578 967
rect 19904 960 20455 967
rect 23681 960 23973 967
rect 14392 926 19578 960
rect 14392 874 14430 926
rect 14482 874 14641 926
rect 14693 874 14852 926
rect 14904 923 18434 926
rect 14904 877 15215 923
rect 15261 877 15373 923
rect 15419 877 15531 923
rect 15577 877 15689 923
rect 15735 877 15847 923
rect 15893 877 16005 923
rect 16051 877 16164 923
rect 16210 877 16322 923
rect 16368 877 16480 923
rect 16526 877 16638 923
rect 16684 877 16796 923
rect 16842 877 16954 923
rect 17000 877 17112 923
rect 17158 877 17271 923
rect 17317 877 17429 923
rect 17475 877 17587 923
rect 17633 877 17745 923
rect 17791 877 17903 923
rect 17949 877 18061 923
rect 18107 877 18434 923
rect 14904 874 18434 877
rect 18486 874 18644 926
rect 18696 874 18855 926
rect 18907 874 19067 926
rect 19119 874 19278 926
rect 19330 874 19488 926
rect 19540 874 19578 926
rect 14392 840 19578 874
rect 19903 926 20455 960
rect 19903 874 19942 926
rect 19994 874 20153 926
rect 20205 874 20364 926
rect 20416 874 20455 926
rect 19903 840 20455 874
rect 23479 840 23973 960
rect 14392 833 14942 840
rect 12958 782 13120 793
rect 9333 688 9462 728
rect 9333 636 9371 688
rect 9423 636 9462 688
rect 9333 609 9462 636
rect 9842 710 9958 747
rect 12958 736 12969 782
rect 13109 736 13120 782
rect 12958 729 13120 736
rect 9842 664 9877 710
rect 9923 664 9958 710
rect 9333 596 9461 609
rect 9519 473 9681 513
rect 9519 421 9590 473
rect 9642 421 9681 473
rect 7449 198 7757 203
rect 6034 78 6549 198
rect 7035 162 7757 198
rect 7035 110 7487 162
rect 7539 110 7667 162
rect 7719 110 7757 162
rect 7035 78 7757 110
rect 7449 70 7757 78
rect 8254 178 8322 300
rect 9519 290 9681 421
rect 9405 287 9681 290
rect 9405 279 9590 287
rect 9405 233 9440 279
rect 9486 235 9590 279
rect 9642 266 9681 287
rect 9842 266 9958 664
rect 10314 595 13120 729
rect 15180 759 18142 840
rect 18396 833 19578 840
rect 19904 833 20455 840
rect 15180 713 15215 759
rect 15261 713 15373 759
rect 15419 713 15531 759
rect 15577 713 15689 759
rect 15735 713 15847 759
rect 15893 713 16005 759
rect 16051 713 16164 759
rect 16210 713 16322 759
rect 16368 713 16480 759
rect 16526 713 16638 759
rect 16684 713 16796 759
rect 16842 713 16954 759
rect 17000 713 17112 759
rect 17158 713 17271 759
rect 17317 713 17429 759
rect 17475 713 17587 759
rect 17633 713 17745 759
rect 17791 713 17903 759
rect 17949 713 18061 759
rect 18107 713 18142 759
rect 23681 799 23973 840
rect 23681 753 23819 799
rect 23865 753 23973 799
rect 14201 653 14466 699
rect 15180 677 18142 713
rect 20631 702 20939 743
rect 13937 587 14105 598
rect 13937 541 13954 587
rect 14094 541 14105 587
rect 13937 497 14105 541
rect 11825 364 14105 497
rect 14201 266 14317 653
rect 18501 627 19473 667
rect 18501 575 18539 627
rect 18591 575 18750 627
rect 18802 575 18961 627
rect 19013 575 19172 627
rect 19224 575 19383 627
rect 19435 575 19473 627
rect 20631 650 20669 702
rect 20721 650 20849 702
rect 20901 650 20939 702
rect 20631 610 20939 650
rect 21185 727 21253 738
rect 18153 520 18283 561
rect 18501 535 19473 575
rect 14497 464 14837 504
rect 14497 412 14535 464
rect 14587 412 14747 464
rect 14799 412 14837 464
rect 14497 371 14837 412
rect 18153 468 18192 520
rect 18244 468 18283 520
rect 18153 465 18283 468
rect 14996 356 17975 389
rect 14996 310 15060 356
rect 15200 310 17975 356
rect 9642 235 14514 266
rect 14996 255 17975 310
rect 18153 325 18218 465
rect 18264 325 18283 465
rect 19858 464 20408 504
rect 18153 302 18283 325
rect 19416 310 19756 429
rect 19858 412 19896 464
rect 19948 412 20107 464
rect 20159 412 20318 464
rect 20370 412 20408 464
rect 19858 371 20408 412
rect 9486 233 14514 235
rect 9405 230 14514 233
rect 9405 184 13335 230
rect 13381 184 13502 230
rect 13548 184 13667 230
rect 13713 184 13832 230
rect 13878 184 14514 230
rect 18153 250 18192 302
rect 18244 250 18283 302
rect 18153 210 18283 250
rect 19640 253 19756 310
rect 21185 305 21196 727
rect 21242 305 21253 727
rect 21393 695 21701 736
rect 21393 643 21431 695
rect 21483 643 21611 695
rect 21663 643 21701 695
rect 21393 603 21701 643
rect 23681 635 23973 753
rect 23681 589 23819 635
rect 23865 589 23973 635
rect 23681 497 23973 589
rect 23181 378 23973 497
rect 21185 253 21253 305
rect 19640 216 21253 253
rect 4313 26 4621 67
rect 8254 58 9319 178
rect 9405 146 14514 184
rect 18501 164 19473 204
rect 18501 112 18539 164
rect 18591 112 18750 164
rect 18802 112 18961 164
rect 19013 112 19172 164
rect 19224 112 19383 164
rect 19435 112 19473 164
rect 19640 170 20112 216
rect 20158 170 20299 216
rect 20345 170 20486 216
rect 20532 170 20672 216
rect 20718 170 20859 216
rect 20905 170 21253 216
rect 19640 160 21253 170
rect 20077 133 21253 160
rect 21393 232 21701 273
rect 21393 180 21431 232
rect 21483 180 21611 232
rect 21663 180 21701 232
rect 21393 140 21701 180
rect 23681 146 23973 378
rect 18501 72 19473 112
rect 23681 100 23819 146
rect 23865 100 23973 146
rect 19695 67 19851 74
rect 4313 -26 4351 26
rect 4403 23 4531 26
rect 4403 -23 4512 23
rect 4403 -26 4531 -23
rect 4583 -26 4621 26
rect 4313 -66 4621 -26
rect 4466 -74 4621 -66
rect 19695 26 20004 67
rect 19695 -26 19734 26
rect 19786 23 19914 26
rect 19802 -23 19914 23
rect 19786 -26 19914 -23
rect 19966 -26 20004 26
rect 19695 -66 20004 -26
rect 19695 -74 19851 -66
rect 23681 -67 23973 100
<< via1 >>
rect 3880 874 3932 926
rect 4091 874 4143 926
rect 4303 874 4355 926
rect 4514 874 4566 926
rect 4816 874 4868 926
rect 5026 874 5078 926
rect 5237 874 5289 926
rect 5449 874 5501 926
rect 5660 874 5712 926
rect 5870 874 5922 926
rect 7926 923 7978 926
rect 7926 877 7978 923
rect 7926 874 7978 877
rect 8137 874 8189 926
rect 8348 874 8400 926
rect 8648 923 8700 926
rect 8828 923 8880 926
rect 8648 877 8658 923
rect 8658 877 8700 923
rect 8828 877 8862 923
rect 8862 877 8880 923
rect 8648 874 8700 877
rect 8828 874 8880 877
rect 2653 650 2705 702
rect 2833 650 2885 702
rect 3415 658 3467 710
rect 3595 658 3647 710
rect 4928 572 4980 624
rect 5139 572 5191 624
rect 5350 572 5402 624
rect 5561 572 5613 624
rect 5772 572 5824 624
rect 7487 584 7539 636
rect 7667 584 7719 636
rect 3863 412 3915 464
rect 4043 412 4095 464
rect 4223 412 4275 464
rect 2653 202 2705 254
rect 2833 202 2885 254
rect 4928 112 4980 164
rect 5139 112 5191 164
rect 5350 112 5402 164
rect 5561 112 5613 164
rect 5772 112 5824 164
rect 6274 337 6293 389
rect 6293 337 6326 389
rect 6557 344 6609 396
rect 6768 344 6820 396
rect 6980 344 7032 396
rect 7191 344 7243 396
rect 9849 874 9901 926
rect 10029 874 10081 926
rect 13386 874 13438 926
rect 13597 874 13649 926
rect 13809 923 13861 926
rect 13809 877 13832 923
rect 13832 877 13861 923
rect 13809 874 13861 877
rect 14020 874 14072 926
rect 14430 874 14482 926
rect 14641 874 14693 926
rect 14852 874 14904 926
rect 18434 874 18486 926
rect 18644 874 18696 926
rect 18855 874 18907 926
rect 19067 874 19119 926
rect 19278 874 19330 926
rect 19488 874 19540 926
rect 19942 874 19994 926
rect 20153 874 20205 926
rect 20364 874 20416 926
rect 9371 636 9423 688
rect 9590 421 9642 473
rect 7487 110 7539 162
rect 7667 110 7719 162
rect 9590 235 9642 287
rect 18539 575 18591 627
rect 18750 575 18802 627
rect 18961 575 19013 627
rect 19172 575 19224 627
rect 19383 575 19435 627
rect 20669 650 20721 702
rect 20849 650 20901 702
rect 14535 412 14587 464
rect 14747 412 14799 464
rect 18192 468 18244 520
rect 19896 412 19948 464
rect 20107 412 20159 464
rect 20318 412 20370 464
rect 18192 250 18244 302
rect 21431 643 21483 695
rect 21611 643 21663 695
rect 18539 112 18591 164
rect 18750 112 18802 164
rect 18961 112 19013 164
rect 19172 112 19224 164
rect 19383 112 19435 164
rect 21431 180 21483 232
rect 21611 180 21663 232
rect 4351 -26 4403 26
rect 4531 23 4583 26
rect 4531 -23 4558 23
rect 4558 -23 4583 23
rect 4531 -26 4583 -23
rect 19734 23 19786 26
rect 19734 -23 19756 23
rect 19756 -23 19786 23
rect 19734 -26 19786 -23
rect 19914 -26 19966 26
<< metal2 >>
rect 366 -101 2485 1051
rect 3824 926 4621 1051
rect 3824 874 3880 926
rect 3932 874 4091 926
rect 4143 874 4303 926
rect 4355 874 4514 926
rect 4566 874 4621 926
rect 2615 702 2923 743
rect 2615 650 2653 702
rect 2705 650 2833 702
rect 2885 650 2923 702
rect 2615 495 2923 650
rect 2615 439 2651 495
rect 2707 439 2831 495
rect 2887 439 2923 495
rect 2615 254 2923 439
rect 3327 710 3686 751
rect 3327 658 3415 710
rect 3467 658 3595 710
rect 3647 658 3686 710
rect 3327 488 3686 658
rect 3327 432 3413 488
rect 3469 432 3593 488
rect 3649 432 3686 488
rect 3327 359 3686 432
rect 3824 464 4621 874
rect 3824 412 3863 464
rect 3915 412 4043 464
rect 4095 412 4223 464
rect 4275 412 4621 464
rect 2615 202 2653 254
rect 2705 202 2833 254
rect 2885 202 2923 254
rect 2615 162 2923 202
rect 3824 28 4621 412
rect 3824 -28 3878 28
rect 3934 -28 4089 28
rect 4145 -28 4301 28
rect 4357 26 4512 28
rect 4568 26 4621 28
rect 4403 -26 4512 26
rect 4583 -26 4621 26
rect 4357 -28 4512 -26
rect 4568 -28 4621 -26
rect 3824 -101 4621 -28
rect 4727 928 6011 1051
rect 4727 872 4814 928
rect 4870 872 5024 928
rect 5080 872 5235 928
rect 5291 872 5447 928
rect 5503 872 5658 928
rect 5714 872 5868 928
rect 5924 872 6011 928
rect 4727 624 6011 872
rect 4727 572 4928 624
rect 4980 572 5139 624
rect 5191 572 5350 624
rect 5402 572 5561 624
rect 5613 572 5772 624
rect 5824 572 6011 624
rect 4727 164 6011 572
rect 6236 536 6364 575
rect 6236 480 6272 536
rect 6328 513 6364 536
rect 6328 480 6365 513
rect 6236 389 6365 480
rect 6236 337 6274 389
rect 6326 337 6365 389
rect 6236 296 6365 337
rect 6460 396 7340 1051
rect 7865 926 8460 1051
rect 7865 874 7926 926
rect 7978 874 8137 926
rect 8189 874 8348 926
rect 8400 874 8460 926
rect 6460 344 6557 396
rect 6609 344 6768 396
rect 6820 344 6980 396
rect 7032 344 7191 396
rect 7243 344 7340 396
rect 4727 112 4928 164
rect 4980 112 5139 164
rect 5191 112 5350 164
rect 5402 112 5561 164
rect 5613 112 5772 164
rect 5824 112 6011 164
rect 4727 -101 6011 112
rect 6460 -101 7340 344
rect 7448 636 7757 677
rect 7448 584 7487 636
rect 7539 584 7667 636
rect 7719 584 7757 636
rect 7448 305 7757 584
rect 7448 249 7485 305
rect 7541 249 7665 305
rect 7721 249 7757 305
rect 7448 162 7757 249
rect 7448 110 7487 162
rect 7539 110 7667 162
rect 7719 110 7757 162
rect 7448 69 7757 110
rect 7865 28 8460 874
rect 7865 -28 7924 28
rect 7980 -28 8135 28
rect 8191 -28 8346 28
rect 8402 -28 8460 28
rect 7865 -101 8460 -28
rect 8563 928 9215 1051
rect 8563 872 8646 928
rect 8702 872 8826 928
rect 8882 872 9215 928
rect 8563 -101 9215 872
rect 9811 926 10120 1051
rect 9811 874 9849 926
rect 9901 874 10029 926
rect 10081 874 10120 926
rect 9332 688 9461 729
rect 9332 636 9371 688
rect 9423 636 9461 688
rect 9332 305 9461 636
rect 9332 249 9369 305
rect 9425 249 9461 305
rect 9332 210 9461 249
rect 9552 536 9680 575
rect 9552 480 9588 536
rect 9644 514 9680 536
rect 9644 480 9681 514
rect 9552 473 9681 480
rect 9552 421 9590 473
rect 9642 421 9681 473
rect 9552 287 9681 421
rect 9552 235 9590 287
rect 9642 235 9681 287
rect 9552 194 9681 235
rect 9811 28 10120 874
rect 9811 -28 9847 28
rect 9903 -28 10027 28
rect 10083 -28 10120 28
rect 9811 -101 10120 -28
rect 10314 -223 10535 1051
rect 10691 -223 10913 1051
rect 11069 -223 11291 1064
rect 11447 -223 11668 1064
rect 11825 -223 12046 1064
rect 12202 -223 12424 1064
rect 12580 -223 12801 1064
rect 12958 -223 13179 1064
rect 13300 926 14159 1051
rect 13300 874 13386 926
rect 13438 874 13597 926
rect 13649 874 13809 926
rect 13861 874 14020 926
rect 14072 874 14159 926
rect 13300 28 14159 874
rect 13300 -28 13384 28
rect 13440 -28 13595 28
rect 13651 -28 13807 28
rect 13863 -28 14018 28
rect 14074 -28 14159 28
rect 13300 -205 14159 -28
rect 14354 928 14980 1051
rect 14354 872 14428 928
rect 14484 872 14639 928
rect 14695 872 14850 928
rect 14906 872 14980 928
rect 14354 464 14980 872
rect 14354 412 14535 464
rect 14587 412 14747 464
rect 14799 412 14980 464
rect 14354 -205 14980 412
rect 15110 -223 15331 1064
rect 15487 -223 15709 1064
rect 15865 -223 16087 1064
rect 16243 -223 16464 1064
rect 16621 -223 16842 1064
rect 16998 -223 17220 1064
rect 17376 -223 17598 1064
rect 17754 -223 17975 1064
rect 18386 928 19587 1051
rect 18386 872 18432 928
rect 18488 872 18642 928
rect 18698 872 18853 928
rect 18909 872 19065 928
rect 19121 872 19276 928
rect 19332 872 19486 928
rect 19542 872 19587 928
rect 18386 627 19587 872
rect 18386 575 18539 627
rect 18591 575 18750 627
rect 18802 575 18961 627
rect 19013 575 19172 627
rect 19224 575 19383 627
rect 19435 575 19587 627
rect 18153 522 18283 561
rect 18153 466 18190 522
rect 18246 466 18283 522
rect 18153 304 18283 466
rect 18153 248 18190 304
rect 18246 248 18283 304
rect 18153 210 18283 248
rect 18386 164 19587 575
rect 18386 112 18539 164
rect 18591 112 18750 164
rect 18802 112 18961 164
rect 19013 112 19172 164
rect 19224 112 19383 164
rect 19435 112 19587 164
rect 18386 -101 19587 112
rect 19695 926 20509 1051
rect 19695 874 19942 926
rect 19994 874 20153 926
rect 20205 874 20364 926
rect 20416 874 20509 926
rect 19695 464 20509 874
rect 19695 412 19896 464
rect 19948 412 20107 464
rect 20159 412 20318 464
rect 20370 412 20509 464
rect 19695 28 20509 412
rect 20630 702 20940 743
rect 20630 650 20669 702
rect 20721 650 20849 702
rect 20901 650 20940 702
rect 20630 488 20940 650
rect 20630 432 20667 488
rect 20723 432 20847 488
rect 20903 432 20940 488
rect 20630 359 20940 432
rect 21392 695 21702 736
rect 21392 643 21431 695
rect 21483 643 21611 695
rect 21663 643 21702 695
rect 21392 488 21702 643
rect 21392 432 21429 488
rect 21485 432 21609 488
rect 21665 432 21702 488
rect 21392 232 21702 432
rect 21392 180 21431 232
rect 21483 180 21611 232
rect 21663 180 21702 232
rect 21392 140 21702 180
rect 19695 26 19757 28
rect 19813 26 19968 28
rect 19695 -26 19734 26
rect 19813 -26 19914 26
rect 19966 -26 19968 26
rect 19695 -28 19757 -26
rect 19813 -28 19968 -26
rect 20024 -28 20180 28
rect 20236 -28 20391 28
rect 20447 -28 20509 28
rect 19695 -101 20509 -28
rect 21823 -101 23951 1051
<< via2 >>
rect 2651 439 2707 495
rect 2831 439 2887 495
rect 3413 432 3469 488
rect 3593 432 3649 488
rect 3878 -28 3934 28
rect 4089 -28 4145 28
rect 4301 26 4357 28
rect 4512 26 4568 28
rect 4301 -26 4351 26
rect 4351 -26 4357 26
rect 4512 -26 4531 26
rect 4531 -26 4568 26
rect 4301 -28 4357 -26
rect 4512 -28 4568 -26
rect 4814 926 4870 928
rect 4814 874 4816 926
rect 4816 874 4868 926
rect 4868 874 4870 926
rect 4814 872 4870 874
rect 5024 926 5080 928
rect 5024 874 5026 926
rect 5026 874 5078 926
rect 5078 874 5080 926
rect 5024 872 5080 874
rect 5235 926 5291 928
rect 5235 874 5237 926
rect 5237 874 5289 926
rect 5289 874 5291 926
rect 5235 872 5291 874
rect 5447 926 5503 928
rect 5447 874 5449 926
rect 5449 874 5501 926
rect 5501 874 5503 926
rect 5447 872 5503 874
rect 5658 926 5714 928
rect 5658 874 5660 926
rect 5660 874 5712 926
rect 5712 874 5714 926
rect 5658 872 5714 874
rect 5868 926 5924 928
rect 5868 874 5870 926
rect 5870 874 5922 926
rect 5922 874 5924 926
rect 5868 872 5924 874
rect 6272 480 6328 536
rect 7485 249 7541 305
rect 7665 249 7721 305
rect 7924 -28 7980 28
rect 8135 -28 8191 28
rect 8346 -28 8402 28
rect 8646 926 8702 928
rect 8646 874 8648 926
rect 8648 874 8700 926
rect 8700 874 8702 926
rect 8646 872 8702 874
rect 8826 926 8882 928
rect 8826 874 8828 926
rect 8828 874 8880 926
rect 8880 874 8882 926
rect 8826 872 8882 874
rect 9369 249 9425 305
rect 9588 480 9644 536
rect 9847 -28 9903 28
rect 10027 -28 10083 28
rect 13384 -28 13440 28
rect 13595 -28 13651 28
rect 13807 -28 13863 28
rect 14018 -28 14074 28
rect 14428 926 14484 928
rect 14428 874 14430 926
rect 14430 874 14482 926
rect 14482 874 14484 926
rect 14428 872 14484 874
rect 14639 926 14695 928
rect 14639 874 14641 926
rect 14641 874 14693 926
rect 14693 874 14695 926
rect 14639 872 14695 874
rect 14850 926 14906 928
rect 14850 874 14852 926
rect 14852 874 14904 926
rect 14904 874 14906 926
rect 14850 872 14906 874
rect 18432 926 18488 928
rect 18432 874 18434 926
rect 18434 874 18486 926
rect 18486 874 18488 926
rect 18432 872 18488 874
rect 18642 926 18698 928
rect 18642 874 18644 926
rect 18644 874 18696 926
rect 18696 874 18698 926
rect 18642 872 18698 874
rect 18853 926 18909 928
rect 18853 874 18855 926
rect 18855 874 18907 926
rect 18907 874 18909 926
rect 18853 872 18909 874
rect 19065 926 19121 928
rect 19065 874 19067 926
rect 19067 874 19119 926
rect 19119 874 19121 926
rect 19065 872 19121 874
rect 19276 926 19332 928
rect 19276 874 19278 926
rect 19278 874 19330 926
rect 19330 874 19332 926
rect 19276 872 19332 874
rect 19486 926 19542 928
rect 19486 874 19488 926
rect 19488 874 19540 926
rect 19540 874 19542 926
rect 19486 872 19542 874
rect 18190 520 18246 522
rect 18190 468 18192 520
rect 18192 468 18244 520
rect 18244 468 18246 520
rect 18190 466 18246 468
rect 18190 302 18246 304
rect 18190 250 18192 302
rect 18192 250 18244 302
rect 18244 250 18246 302
rect 18190 248 18246 250
rect 20667 432 20723 488
rect 20847 432 20903 488
rect 21429 432 21485 488
rect 21609 432 21665 488
rect 19757 26 19813 28
rect 19757 -26 19786 26
rect 19786 -26 19813 26
rect 19757 -28 19813 -26
rect 19968 -28 20024 28
rect 20180 -28 20236 28
rect 20391 -28 20447 28
<< metal3 >>
rect -1 928 24218 1001
rect -1 872 4814 928
rect 4870 872 5024 928
rect 5080 872 5235 928
rect 5291 872 5447 928
rect 5503 872 5658 928
rect 5714 872 5868 928
rect 5924 872 8646 928
rect 8702 872 8826 928
rect 8882 872 14428 928
rect 14484 872 14639 928
rect 14695 872 14850 928
rect 14906 872 18432 928
rect 18488 872 18642 928
rect 18698 872 18853 928
rect 18909 872 19065 928
rect 19121 872 19276 928
rect 19332 872 19486 928
rect 19542 872 24218 928
rect -1 799 24218 872
rect 6244 574 9637 575
rect -1 495 3686 561
rect -1 439 2651 495
rect 2707 439 2831 495
rect 2887 488 3686 495
rect 2887 439 3413 488
rect -1 432 3413 439
rect 3469 432 3593 488
rect 3649 432 3686 488
rect 6236 536 9681 574
rect 6236 480 6272 536
rect 6328 480 9588 536
rect 9644 480 9681 536
rect 6236 441 9681 480
rect 18153 522 18283 561
rect 18153 466 18190 522
rect 18246 466 18283 522
rect -1 359 3686 432
rect 18153 343 18283 466
rect 20630 488 24218 561
rect 20630 432 20667 488
rect 20723 432 20847 488
rect 20903 432 21429 488
rect 21485 432 21609 488
rect 21665 432 24218 488
rect 20630 359 24218 432
rect 7448 305 18283 343
rect 7448 249 7485 305
rect 7541 249 7665 305
rect 7721 249 9369 305
rect 9425 304 18283 305
rect 9425 249 18190 304
rect 7448 248 18190 249
rect 18246 248 18283 304
rect 7448 210 18283 248
rect -1 28 24218 101
rect -1 -28 3878 28
rect 3934 -28 4089 28
rect 4145 -28 4301 28
rect 4357 -28 4512 28
rect 4568 -28 7924 28
rect 7980 -28 8135 28
rect 8191 -28 8346 28
rect 8402 -28 9847 28
rect 9903 -28 10027 28
rect 10083 -28 13384 28
rect 13440 -28 13595 28
rect 13651 -28 13807 28
rect 13863 -28 14018 28
rect 14074 -28 19757 28
rect 19813 -28 19968 28
rect 20024 -28 20180 28
rect 20236 -28 20391 28
rect 20447 -28 24218 28
rect -1 -101 24218 -28
use M1_NWELL$$46890028_64x8m81  M1_NWELL$$46890028_64x8m81_0
timestamp 1666464484
transform 1 0 8760 0 1 900
box 0 0 1 1
use M1_NWELL4310589983236_64x8m81  M1_NWELL4310589983236_64x8m81_0
timestamp 1666464484
transform 1 0 6202 0 1 900
box 0 0 1 1
use M1_PACTIVE$$204209196_64x8m81  M1_PACTIVE$$204209196_64x8m81_0
timestamp 1666464484
transform 1 0 4535 0 1 0
box 0 0 1 1
use M1_PACTIVE43105899832103_64x8m81  M1_PACTIVE43105899832103_64x8m81_0
timestamp 1666464484
transform 1 0 7811 0 1 900
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1666464484
transform 1 0 9900 0 1 687
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_1
timestamp 1666464484
transform 1 0 9463 0 1 256
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_0
timestamp 1666464484
transform 1 0 14024 0 1 564
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_1
timestamp 1666464484
transform 1 0 13039 0 1 759
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1666464484
transform 0 1 15130 -1 0 333
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_1
timestamp 1666464484
transform 1 0 6316 0 1 368
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_2
timestamp 1666464484
transform 1 0 8288 0 1 370
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_3
timestamp 1666464484
transform 1 0 18241 0 1 395
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_4
timestamp 1666464484
transform 1 0 6094 0 1 368
box 0 0 1 1
use M1_POLY243105899832102_64x8m81  M1_POLY243105899832102_64x8m81_0
timestamp 1666464484
transform 1 0 21219 0 1 516
box 0 0 1 1
use M1_POLY243105899832102_64x8m81  M1_POLY243105899832102_64x8m81_1
timestamp 1666464484
transform 1 0 3114 0 1 546
box 0 0 1 1
use M1_PSUB$$45111340_64x8m81  M1_PSUB$$45111340_64x8m81_0
timestamp 1666464484
transform -1 0 19779 0 1 0
box 0 0 1 1
use M1_PSUB$$49279020_64x8m81  M1_PSUB$$49279020_64x8m81_0
timestamp 1666464484
transform 1 0 11483 0 1 900
box -1108 -83 1108 83
use M2_M1$$45004844_64x8m81  M2_M1$$45004844_64x8m81_0
timestamp 1666464484
transform 1 0 20179 0 1 900
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_0
timestamp 1666464484
transform 1 0 6300 0 1 363
box 0 0 1 1
use M2_M1$$201262124_64x8m81  M2_M1$$201262124_64x8m81_0
timestamp 1666464484
transform 1 0 14667 0 1 438
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_0
timestamp 1666464484
transform 1 0 6300 0 1 363
box 0 0 1 1
use M2_M1$$202394668_64x8m81  M2_M1$$202394668_64x8m81_1
timestamp 1666464484
transform 1 0 9397 0 1 662
box 0 0 1 1
use M2_M1$$202406956_64x8m81  M2_M1$$202406956_64x8m81_0
timestamp 1666464484
transform 1 0 18218 0 1 385
box 0 0 1 1
use M2_M1$$204402732_64x8m81  M2_M1$$204402732_64x8m81_0
timestamp 1666464484
transform 1 0 22887 0 1 0
box -1013 -67 1013 67
use M2_M1$$204402732_64x8m81  M2_M1$$204402732_64x8m81_1
timestamp 1666464484
transform 1 0 22887 0 1 900
box -1013 -67 1013 67
use M2_M1$$204402732_64x8m81  M2_M1$$204402732_64x8m81_2
timestamp 1666464484
transform 1 0 1425 0 1 0
box -1013 -67 1013 67
use M2_M1$$204402732_64x8m81  M2_M1$$204402732_64x8m81_3
timestamp 1666464484
transform 1 0 1425 0 1 900
box -1013 -67 1013 67
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_0
timestamp 1666464484
transform 1 0 7603 0 1 610
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_1
timestamp 1666464484
transform 1 0 9965 0 1 900
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_2
timestamp 1666464484
transform 1 0 21547 0 1 669
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_3
timestamp 1666464484
transform 1 0 19850 0 1 0
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_4
timestamp 1666464484
transform 1 0 8764 0 1 900
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_5
timestamp 1666464484
transform 1 0 4467 0 1 0
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_6
timestamp 1666464484
transform 1 0 7603 0 1 136
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_7
timestamp 1666464484
transform 1 0 20785 0 1 676
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_8
timestamp 1666464484
transform 1 0 2769 0 1 676
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_9
timestamp 1666464484
transform 1 0 2769 0 1 228
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_10
timestamp 1666464484
transform 1 0 3531 0 1 684
box 0 0 1 1
use M2_M1$$204403756_64x8m81  M2_M1$$204403756_64x8m81_11
timestamp 1666464484
transform 1 0 21547 0 1 206
box 0 0 1 1
use M2_M1$$204403756_R270_64x8m81  M2_M1$$204403756_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 9616 1 0 354
box 0 0 1 1
use M2_M1$$204404780_64x8m81  M2_M1$$204404780_64x8m81_0
timestamp 1666464484
transform 1 0 13729 0 1 900
box 0 0 1 1
use M2_M1$$204404780_64x8m81  M2_M1$$204404780_64x8m81_1
timestamp 1666464484
transform 1 0 4223 0 1 900
box 0 0 1 1
use M2_M1$$204404780_64x8m81  M2_M1$$204404780_64x8m81_2
timestamp 1666464484
transform 1 0 6900 0 1 370
box 0 0 1 1
use M2_M1$$204405804_64x8m81  M2_M1$$204405804_64x8m81_0
timestamp 1666464484
transform 1 0 4069 0 1 438
box 0 0 1 1
use M2_M1$$204406828_64x8m81  M2_M1$$204406828_64x8m81_0
timestamp 1666464484
transform 1 0 18987 0 1 900
box 0 0 1 1
use M2_M1$$204406828_64x8m81  M2_M1$$204406828_64x8m81_1
timestamp 1666464484
transform 1 0 5369 0 1 900
box 0 0 1 1
use M2_M1$$204407852_64x8m81  M2_M1$$204407852_64x8m81_0
timestamp 1666464484
transform 1 0 5376 0 1 598
box 0 0 1 1
use M2_M1$$204407852_64x8m81  M2_M1$$204407852_64x8m81_1
timestamp 1666464484
transform 1 0 5376 0 1 138
box 0 0 1 1
use M2_M1$$204407852_64x8m81  M2_M1$$204407852_64x8m81_2
timestamp 1666464484
transform 1 0 18987 0 1 601
box 0 0 1 1
use M2_M1$$204407852_64x8m81  M2_M1$$204407852_64x8m81_3
timestamp 1666464484
transform 1 0 18987 0 1 138
box 0 0 1 1
use M2_M1$$204408876_64x8m81  M2_M1$$204408876_64x8m81_0
timestamp 1666464484
transform 1 0 14667 0 1 900
box 0 0 1 1
use M2_M1$$204408876_64x8m81  M2_M1$$204408876_64x8m81_1
timestamp 1666464484
transform 1 0 20133 0 1 438
box 0 0 1 1
use M2_M1$$204408876_64x8m81  M2_M1$$204408876_64x8m81_2
timestamp 1666464484
transform 1 0 8163 0 1 900
box 0 0 1 1
use M3_M2$$201251884_64x8m81  M3_M2$$201251884_64x8m81_0
timestamp 1666464484
transform 1 0 20102 0 1 0
box 0 0 1 1
use M3_M2$$201251884_64x8m81  M3_M2$$201251884_64x8m81_1
timestamp 1666464484
transform 1 0 13729 0 1 0
box 0 0 1 1
use M3_M2$$201251884_64x8m81  M3_M2$$201251884_64x8m81_2
timestamp 1666464484
transform 1 0 4223 0 1 0
box 0 0 1 1
use M3_M2$$201252908_64x8m81  M3_M2$$201252908_64x8m81_0
timestamp 1666464484
transform 1 0 18218 0 1 385
box 0 0 1 1
use M3_M2$$204147756_64x8m81  M3_M2$$204147756_64x8m81_0
timestamp 1666464484
transform 1 0 14667 0 1 900
box 0 0 1 1
use M3_M2$$204147756_64x8m81  M3_M2$$204147756_64x8m81_1
timestamp 1666464484
transform 1 0 8163 0 1 0
box 0 0 1 1
use M3_M2$$204398636_64x8m81  M3_M2$$204398636_64x8m81_0
timestamp 1666464484
transform 1 0 9616 0 1 508
box 0 0 1 1
use M3_M2$$204398636_64x8m81  M3_M2$$204398636_64x8m81_1
timestamp 1666464484
transform 1 0 6300 0 1 508
box 0 0 1 1
use M3_M2$$204398636_64x8m81  M3_M2$$204398636_64x8m81_2
timestamp 1666464484
transform 1 0 9397 0 1 277
box 0 0 1 1
use M3_M2$$204399660_64x8m81  M3_M2$$204399660_64x8m81_0
timestamp 1666464484
transform 1 0 22887 0 1 900
box -1013 -67 1013 67
use M3_M2$$204399660_64x8m81  M3_M2$$204399660_64x8m81_1
timestamp 1666464484
transform 1 0 1425 0 1 900
box -1013 -67 1013 67
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_0
timestamp 1666464484
transform 1 0 9965 0 1 0
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_1
timestamp 1666464484
transform 1 0 7603 0 1 277
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_2
timestamp 1666464484
transform 1 0 2769 0 1 467
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_3
timestamp 1666464484
transform 1 0 3531 0 1 460
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_4
timestamp 1666464484
transform 1 0 20785 0 1 460
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_5
timestamp 1666464484
transform 1 0 8764 0 1 900
box 0 0 1 1
use M3_M2$$204400684_64x8m81  M3_M2$$204400684_64x8m81_6
timestamp 1666464484
transform 1 0 21547 0 1 460
box 0 0 1 1
use M3_M2$$204401708_64x8m81  M3_M2$$204401708_64x8m81_0
timestamp 1666464484
transform 1 0 18987 0 1 900
box 0 0 1 1
use M3_M2$$204401708_64x8m81  M3_M2$$204401708_64x8m81_1
timestamp 1666464484
transform 1 0 5369 0 1 900
box 0 0 1 1
use nmos_1p2$$49277996_R270_64x8m81  nmos_1p2$$49277996_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 9763 1 0 759
box -119 -71 177 510
use nmos_5p043105899832107_64x8m81  nmos_5p043105899832107_64x8m81_0
timestamp 1666464484
transform 0 -1 9326 1 0 193
box -88 -44 208 176
use nmos_5p043105899832109_64x8m81  nmos_5p043105899832109_64x8m81_0
timestamp 1666464484
transform 0 -1 4267 -1 0 848
box -88 -44 432 1044
use nmos_5p043105899832109_64x8m81  nmos_5p043105899832109_64x8m81_1
timestamp 1666464484
transform 0 1 20050 -1 0 848
box -88 -44 432 1044
use nmos_5p043105899832110_64x8m81  nmos_5p043105899832110_64x8m81_0
timestamp 1666464484
transform 0 -1 8152 1 0 193
box -88 -44 432 704
use pmos_1p2$$49270828_R270_64x8m81  pmos_1p2$$49270828_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 2932 1 0 311
box -296 -137 817 2333
use pmos_1p2$$49271852_R270_64x8m81  pmos_1p2$$49271852_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 7097 1 0 224
box -296 -137 853 796
use pmos_1p2$$49272876_R270_64x8m81  pmos_1p2$$49272876_R270_64x8m81_0
timestamp 1666464484
transform 0 1 18361 1 0 224
box -296 -137 853 1235
use pmos_1p2$$49272876_R270_64x8m81  pmos_1p2$$49272876_R270_64x8m81_1
timestamp 1666464484
transform 0 -1 5956 1 0 224
box -296 -137 853 1235
use pmos_5p043105899832104_64x8m81  pmos_5p043105899832104_64x8m81_0
timestamp 1666464484
transform 0 1 14395 1 0 504
box -208 -120 328 644
use pmos_5p043105899832104_64x8m81  pmos_5p043105899832104_64x8m81_1
timestamp 1666464484
transform 0 1 14395 1 0 728
box -208 -120 328 644
use pmos_5p043105899832104_64x8m81  pmos_5p043105899832104_64x8m81_2
timestamp 1666464484
transform 0 1 14395 1 0 280
box -208 -120 328 644
use pmos_5p043105899832108_64x8m81  pmos_5p043105899832108_64x8m81_0
timestamp 1666464484
transform 0 1 21385 1 0 280
box -208 -120 776 2120
use pmos_5p043105899832111_64x8m81  pmos_5p043105899832111_64x8m81_0
timestamp 1666464484
transform 0 -1 8922 1 0 193
box -208 -120 328 438
<< labels >>
rlabel metal1 s 13062 662 13062 662 4 xc
port 1 nsew
rlabel metal1 s 13062 431 13062 431 4 xb
port 2 nsew
rlabel metal1 s 15060 322 15060 322 4 xa
port 3 nsew
rlabel metal3 s 195 0 195 0 4 vss
port 4 nsew
rlabel metal3 s 195 900 195 900 4 vdd
port 5 nsew
rlabel metal3 s 23423 460 23423 460 4 RWL
port 6 nsew
rlabel metal3 s 830 460 830 460 4 LWL
port 7 nsew
rlabel metal2 s 6900 855 6900 855 4 men
port 8 nsew
<< properties >>
string GDS_END 1032414
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1015358
<< end >>
