magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -174 44 174 50
rect -174 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 174 44
rect -174 -18 174 18
rect -174 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 174 -18
rect -174 -50 174 -44
<< via1 >>
rect -168 18 -142 44
rect -106 18 -80 44
rect -44 18 -18 44
rect 18 18 44 44
rect 80 18 106 44
rect 142 18 168 44
rect -168 -44 -142 -18
rect -106 -44 -80 -18
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect 80 -44 106 -18
rect 142 -44 168 -18
<< metal2 >>
rect -174 44 174 50
rect -174 18 -168 44
rect -142 18 -106 44
rect -80 18 -44 44
rect -18 18 18 44
rect 44 18 80 44
rect 106 18 142 44
rect 168 18 174 44
rect -174 -18 174 18
rect -174 -44 -168 -18
rect -142 -44 -106 -18
rect -80 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 80 -18
rect 106 -44 142 -18
rect 168 -44 174 -18
rect -174 -50 174 -44
<< properties >>
string GDS_END 1632638
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1631738
<< end >>
