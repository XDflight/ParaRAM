magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -143 169 143 174
rect -143 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 143 169
rect -143 107 143 141
rect -143 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 143 107
rect -143 45 143 79
rect -143 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 143 45
rect -143 -17 143 17
rect -143 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 143 -17
rect -143 -79 143 -45
rect -143 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 143 -79
rect -143 -141 143 -107
rect -143 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 143 -141
rect -143 -174 143 -169
<< via2 >>
rect -138 141 -110 169
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect 110 141 138 169
rect -138 79 -110 107
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect 110 79 138 107
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
rect -138 -107 -110 -79
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect 110 -107 138 -79
rect -138 -169 -110 -141
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect 110 -169 138 -141
<< metal3 >>
rect -143 169 143 174
rect -143 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 143 169
rect -143 107 143 141
rect -143 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 143 107
rect -143 45 143 79
rect -143 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 143 45
rect -143 -17 143 17
rect -143 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 143 -17
rect -143 -79 143 -45
rect -143 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 143 -79
rect -143 -141 143 -107
rect -143 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 143 -141
rect -143 -174 143 -169
<< properties >>
string GDS_END 1802456
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1800404
<< end >>
