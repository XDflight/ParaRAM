magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -170 1007 170 1046
rect -170 951 -134 1007
rect -78 951 78 1007
rect 134 951 170 1007
rect -170 790 170 951
rect -170 734 -134 790
rect -78 734 78 790
rect 134 734 170 790
rect -170 572 170 734
rect -170 516 -134 572
rect -78 516 78 572
rect 134 516 170 572
rect -170 355 170 516
rect -170 299 -134 355
rect -78 299 78 355
rect 134 299 170 355
rect -170 137 170 299
rect -170 81 -134 137
rect -78 81 78 137
rect 134 81 170 137
rect -170 -81 170 81
rect -170 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 170 -81
rect -170 -299 170 -137
rect -170 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 170 -299
rect -170 -516 170 -355
rect -170 -572 -134 -516
rect -78 -572 78 -516
rect 134 -572 170 -516
rect -170 -734 170 -572
rect -170 -790 -134 -734
rect -78 -790 78 -734
rect 134 -790 170 -734
rect -170 -951 170 -790
rect -170 -1007 -134 -951
rect -78 -1007 78 -951
rect 134 -1007 170 -951
rect -170 -1046 170 -1007
<< via2 >>
rect -134 951 -78 1007
rect 78 951 134 1007
rect -134 734 -78 790
rect 78 734 134 790
rect -134 516 -78 572
rect 78 516 134 572
rect -134 299 -78 355
rect 78 299 134 355
rect -134 81 -78 137
rect 78 81 134 137
rect -134 -137 -78 -81
rect 78 -137 134 -81
rect -134 -355 -78 -299
rect 78 -355 134 -299
rect -134 -572 -78 -516
rect 78 -572 134 -516
rect -134 -790 -78 -734
rect 78 -790 134 -734
rect -134 -1007 -78 -951
rect 78 -1007 134 -951
<< metal3 >>
rect -170 1007 170 1046
rect -170 951 -134 1007
rect -78 951 78 1007
rect 134 951 170 1007
rect -170 790 170 951
rect -170 734 -134 790
rect -78 734 78 790
rect 134 734 170 790
rect -170 572 170 734
rect -170 516 -134 572
rect -78 516 78 572
rect 134 516 170 572
rect -170 355 170 516
rect -170 299 -134 355
rect -78 299 78 355
rect 134 299 170 355
rect -170 137 170 299
rect -170 81 -134 137
rect -78 81 78 137
rect 134 81 170 137
rect -170 -81 170 81
rect -170 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 170 -81
rect -170 -299 170 -137
rect -170 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 170 -299
rect -170 -516 170 -355
rect -170 -572 -134 -516
rect -78 -572 78 -516
rect 134 -572 170 -516
rect -170 -734 170 -572
rect -170 -790 -134 -734
rect -78 -790 78 -734
rect 134 -790 170 -734
rect -170 -951 170 -790
rect -170 -1007 -134 -951
rect -78 -1007 78 -951
rect 134 -1007 170 -951
rect -170 -1046 170 -1007
<< properties >>
string GDS_END 684294
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 682882
<< end >>
