magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 51823 242 51842
rect -42 -23 -23 51823
rect 223 -23 242 51823
rect -42 -42 242 -23
<< psubdiffcont >>
rect -23 -23 223 51823
<< metal1 >>
rect -34 51823 234 51834
rect -34 -23 -23 51823
rect 223 -23 234 51823
rect -34 -34 234 -23
<< properties >>
string GDS_END 2036572
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1936728
<< end >>
