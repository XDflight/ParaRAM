magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1990 1094
<< pwell >>
rect -86 -86 1990 453
<< mvnmos >>
rect 124 215 244 333
rect 397 215 517 333
rect 621 215 741 333
rect 997 69 1117 333
rect 1368 215 1488 333
rect 1660 215 1780 333
<< mvpmos >>
rect 124 683 224 881
rect 328 683 428 881
rect 542 683 642 881
rect 1007 576 1107 936
rect 1388 662 1488 860
rect 1660 662 1760 860
<< mvndiff >>
rect 36 285 124 333
rect 36 239 49 285
rect 95 239 124 285
rect 36 215 124 239
rect 244 285 397 333
rect 244 239 322 285
rect 368 239 397 285
rect 244 215 397 239
rect 517 285 621 333
rect 517 239 546 285
rect 592 239 621 285
rect 517 215 621 239
rect 741 285 829 333
rect 741 239 770 285
rect 816 239 829 285
rect 741 215 829 239
rect 909 285 997 333
rect 909 239 922 285
rect 968 239 997 285
rect 909 69 997 239
rect 1117 222 1205 333
rect 1117 82 1146 222
rect 1192 82 1205 222
rect 1280 285 1368 333
rect 1280 239 1293 285
rect 1339 239 1368 285
rect 1280 215 1368 239
rect 1488 285 1660 333
rect 1488 239 1517 285
rect 1563 239 1660 285
rect 1488 215 1660 239
rect 1780 285 1868 333
rect 1780 239 1809 285
rect 1855 239 1868 285
rect 1780 215 1868 239
rect 1117 69 1205 82
<< mvpdiff >>
rect 36 847 124 881
rect 36 707 49 847
rect 95 707 124 847
rect 36 683 124 707
rect 224 847 328 881
rect 224 707 253 847
rect 299 707 328 847
rect 224 683 328 707
rect 428 847 542 881
rect 428 707 467 847
rect 513 707 542 847
rect 428 683 542 707
rect 642 753 730 881
rect 642 707 671 753
rect 717 707 730 753
rect 642 683 730 707
rect 919 769 1007 936
rect 919 629 932 769
rect 978 629 1007 769
rect 919 576 1007 629
rect 1107 923 1195 936
rect 1107 783 1136 923
rect 1182 783 1195 923
rect 1107 576 1195 783
rect 1300 847 1388 860
rect 1300 707 1313 847
rect 1359 707 1388 847
rect 1300 662 1388 707
rect 1488 847 1660 860
rect 1488 707 1517 847
rect 1563 707 1660 847
rect 1488 662 1660 707
rect 1760 847 1848 860
rect 1760 707 1789 847
rect 1835 707 1848 847
rect 1760 662 1848 707
<< mvndiffc >>
rect 49 239 95 285
rect 322 239 368 285
rect 546 239 592 285
rect 770 239 816 285
rect 922 239 968 285
rect 1146 82 1192 222
rect 1293 239 1339 285
rect 1517 239 1563 285
rect 1809 239 1855 285
<< mvpdiffc >>
rect 49 707 95 847
rect 253 707 299 847
rect 467 707 513 847
rect 671 707 717 753
rect 932 629 978 769
rect 1136 783 1182 923
rect 1313 707 1359 847
rect 1517 707 1563 847
rect 1789 707 1835 847
<< polysilicon >>
rect 1007 936 1107 980
rect 124 881 224 925
rect 328 881 428 925
rect 542 881 642 925
rect 124 550 224 683
rect 328 550 428 683
rect 542 650 642 683
rect 542 604 555 650
rect 601 604 642 650
rect 542 591 642 604
rect 1388 860 1488 904
rect 1660 860 1760 904
rect 124 543 517 550
rect 1007 543 1107 576
rect 124 510 741 543
rect 124 449 244 510
rect 494 503 741 510
rect 124 403 137 449
rect 183 403 244 449
rect 124 333 244 403
rect 397 449 469 462
rect 397 403 410 449
rect 456 403 469 449
rect 557 404 741 503
rect 1007 497 1037 543
rect 1083 497 1107 543
rect 1007 484 1107 497
rect 1388 449 1488 662
rect 397 377 469 403
rect 397 333 517 377
rect 621 333 741 404
rect 997 423 1117 436
rect 997 377 1029 423
rect 1075 377 1117 423
rect 1388 403 1429 449
rect 1475 403 1488 449
rect 1388 377 1488 403
rect 997 333 1117 377
rect 1368 333 1488 377
rect 1660 449 1760 662
rect 1660 403 1701 449
rect 1747 403 1760 449
rect 1660 377 1760 403
rect 1660 333 1780 377
rect 124 171 244 215
rect 397 171 517 215
rect 621 171 741 215
rect 1368 171 1488 215
rect 1660 171 1780 215
rect 997 25 1117 69
<< polycontact >>
rect 555 604 601 650
rect 137 403 183 449
rect 410 403 456 449
rect 1037 497 1083 543
rect 1029 377 1075 423
rect 1429 403 1475 449
rect 1701 403 1747 449
<< metal1 >>
rect 0 923 1904 1098
rect 0 918 1136 923
rect 49 847 95 858
rect 49 650 95 707
rect 253 847 299 918
rect 253 696 299 707
rect 467 847 1070 872
rect 513 826 1070 847
rect 467 696 513 707
rect 671 753 717 764
rect 49 604 555 650
rect 601 604 612 650
rect 30 449 194 542
rect 421 449 467 604
rect 30 403 137 449
rect 183 403 194 449
rect 240 403 410 449
rect 456 403 467 449
rect 240 364 286 403
rect 219 325 286 364
rect 219 285 265 325
rect 38 239 49 285
rect 95 239 265 285
rect 322 285 368 296
rect 671 285 717 707
rect 535 239 546 285
rect 592 239 717 285
rect 322 90 368 239
rect 671 182 717 239
rect 770 285 816 826
rect 770 228 816 239
rect 922 769 978 780
rect 922 629 932 769
rect 922 354 978 629
rect 1024 726 1070 826
rect 1182 918 1904 923
rect 1136 772 1182 783
rect 1313 847 1359 858
rect 1024 707 1313 726
rect 1024 680 1359 707
rect 1517 847 1563 918
rect 1517 696 1563 707
rect 1789 847 1835 858
rect 1024 543 1083 680
rect 1789 676 1835 707
rect 1024 497 1037 543
rect 1024 486 1083 497
rect 1609 630 1835 676
rect 1609 449 1655 630
rect 1029 423 1075 434
rect 1418 403 1429 449
rect 1475 403 1655 449
rect 922 285 968 354
rect 1029 325 1075 377
rect 1029 313 1339 325
rect 922 228 968 239
rect 1014 285 1339 313
rect 1014 279 1293 285
rect 1014 182 1060 279
rect 671 136 1060 182
rect 1146 222 1192 233
rect 1293 228 1339 239
rect 1517 285 1563 296
rect 1609 285 1655 403
rect 1701 449 1762 542
rect 1747 403 1762 449
rect 1701 354 1762 403
rect 1609 239 1809 285
rect 1855 239 1866 285
rect 0 82 1146 90
rect 1517 90 1563 239
rect 1192 82 1904 90
rect 0 -90 1904 82
<< labels >>
flabel metal1 s 30 403 194 542 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1701 354 1762 542 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 1904 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 1517 233 1563 296 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 922 354 978 780 0 FreeSans 200 0 0 0 ZN
port 3 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 922 228 968 354 1 ZN
port 3 nsew default output
rlabel metal1 s 1517 772 1563 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1136 772 1182 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 772 299 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1517 696 1563 772 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 253 696 299 772 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 322 233 368 296 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1517 90 1563 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1146 90 1192 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 322 90 368 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1904 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1904 1008
string GDS_END 905838
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 900330
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
