magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -803 26 803 66
rect -803 -26 -764 26
rect -712 -26 -553 26
rect -501 -26 -343 26
rect -291 -26 -132 26
rect -80 -26 80 26
rect 132 -26 291 26
rect 343 -26 501 26
rect 553 -26 712 26
rect 764 -26 803 26
rect -803 -67 803 -26
<< via1 >>
rect -764 -26 -712 26
rect -553 -26 -501 26
rect -343 -26 -291 26
rect -132 -26 -80 26
rect 80 -26 132 26
rect 291 -26 343 26
rect 501 -26 553 26
rect 712 -26 764 26
<< metal2 >>
rect -802 26 803 66
rect -802 -26 -764 26
rect -712 -26 -553 26
rect -501 -26 -343 26
rect -291 -26 -132 26
rect -80 -26 80 26
rect 132 -26 291 26
rect 343 -26 501 26
rect 553 -26 712 26
rect 764 -26 803 26
rect -802 -67 803 -26
<< properties >>
string GDS_END 611096
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 610452
<< end >>
