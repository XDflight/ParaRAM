magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 400
rect 224 0 344 400
rect 448 0 568 400
<< mvndiff >>
rect -88 387 0 400
rect -88 341 -75 387
rect -29 341 0 387
rect -88 278 0 341
rect -88 232 -75 278
rect -29 232 0 278
rect -88 169 0 232
rect -88 123 -75 169
rect -29 123 0 169
rect -88 59 0 123
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 387 224 400
rect 120 341 149 387
rect 195 341 224 387
rect 120 278 224 341
rect 120 232 149 278
rect 195 232 224 278
rect 120 169 224 232
rect 120 123 149 169
rect 195 123 224 169
rect 120 59 224 123
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 387 448 400
rect 344 341 373 387
rect 419 341 448 387
rect 344 278 448 341
rect 344 232 373 278
rect 419 232 448 278
rect 344 169 448 232
rect 344 123 373 169
rect 419 123 448 169
rect 344 59 448 123
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 387 656 400
rect 568 341 597 387
rect 643 341 656 387
rect 568 278 656 341
rect 568 232 597 278
rect 643 232 656 278
rect 568 169 656 232
rect 568 123 597 169
rect 643 123 656 169
rect 568 59 656 123
rect 568 13 597 59
rect 643 13 656 59
rect 568 0 656 13
<< mvndiffc >>
rect -75 341 -29 387
rect -75 232 -29 278
rect -75 123 -29 169
rect -75 13 -29 59
rect 149 341 195 387
rect 149 232 195 278
rect 149 123 195 169
rect 149 13 195 59
rect 373 341 419 387
rect 373 232 419 278
rect 373 123 419 169
rect 373 13 419 59
rect 597 341 643 387
rect 597 232 643 278
rect 597 123 643 169
rect 597 13 643 59
<< polysilicon >>
rect 0 400 120 444
rect 224 400 344 444
rect 448 400 568 444
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
<< metal1 >>
rect -75 387 -29 400
rect -75 278 -29 341
rect -75 169 -29 232
rect -75 59 -29 123
rect -75 0 -29 13
rect 149 387 195 400
rect 149 278 195 341
rect 149 169 195 232
rect 149 59 195 123
rect 149 0 195 13
rect 373 387 419 400
rect 373 278 419 341
rect 373 169 419 232
rect 373 59 419 123
rect 373 0 419 13
rect 597 387 643 400
rect 597 278 643 341
rect 597 169 643 232
rect 597 59 643 123
rect 597 0 643 13
<< labels >>
flabel metal1 s -52 200 -52 200 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 200 620 200 0 FreeSans 200 0 0 0 D
flabel metal1 s 172 200 172 200 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 200 396 200 0 FreeSans 200 0 0 0 S
<< properties >>
string GDS_END 508804
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 506120
<< end >>
