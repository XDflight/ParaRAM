magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1766 1094
<< pwell >>
rect -86 -86 1766 453
<< mvnmos >>
rect 126 69 246 333
rect 350 69 470 333
rect 574 69 694 333
rect 988 68 1108 332
rect 1212 68 1332 332
rect 1436 68 1556 332
<< mvpmos >>
rect 146 573 246 933
rect 350 573 450 933
rect 660 573 760 933
rect 1008 580 1108 940
rect 1212 580 1312 940
rect 1416 580 1516 940
<< mvndiff >>
rect 38 320 126 333
rect 38 180 51 320
rect 97 180 126 320
rect 38 69 126 180
rect 246 222 350 333
rect 246 82 275 222
rect 321 82 350 222
rect 246 69 350 82
rect 470 287 574 333
rect 470 147 499 287
rect 545 147 574 287
rect 470 69 574 147
rect 694 320 782 333
rect 694 274 723 320
rect 769 274 782 320
rect 694 69 782 274
rect 900 206 988 332
rect 900 160 913 206
rect 959 160 988 206
rect 900 68 988 160
rect 1108 221 1212 332
rect 1108 81 1137 221
rect 1183 81 1212 221
rect 1108 68 1212 81
rect 1332 319 1436 332
rect 1332 179 1361 319
rect 1407 179 1436 319
rect 1332 68 1436 179
rect 1556 221 1644 332
rect 1556 81 1585 221
rect 1631 81 1644 221
rect 1556 68 1644 81
<< mvpdiff >>
rect 58 726 146 933
rect 58 586 71 726
rect 117 586 146 726
rect 58 573 146 586
rect 246 920 350 933
rect 246 780 275 920
rect 321 780 350 920
rect 246 573 350 780
rect 450 726 660 933
rect 450 586 585 726
rect 631 586 660 726
rect 450 573 660 586
rect 760 632 848 933
rect 760 586 789 632
rect 835 586 848 632
rect 760 573 848 586
rect 920 639 1008 940
rect 920 593 933 639
rect 979 593 1008 639
rect 920 580 1008 593
rect 1108 927 1212 940
rect 1108 787 1137 927
rect 1183 787 1212 927
rect 1108 580 1212 787
rect 1312 733 1416 940
rect 1312 593 1341 733
rect 1387 593 1416 733
rect 1312 580 1416 593
rect 1516 927 1604 940
rect 1516 787 1545 927
rect 1591 787 1604 927
rect 1516 580 1604 787
<< mvndiffc >>
rect 51 180 97 320
rect 275 82 321 222
rect 499 147 545 287
rect 723 274 769 320
rect 913 160 959 206
rect 1137 81 1183 221
rect 1361 179 1407 319
rect 1585 81 1631 221
<< mvpdiffc >>
rect 71 586 117 726
rect 275 780 321 920
rect 585 586 631 726
rect 789 586 835 632
rect 933 593 979 639
rect 1137 787 1183 927
rect 1341 593 1387 733
rect 1545 787 1591 927
<< polysilicon >>
rect 146 933 246 977
rect 350 933 450 977
rect 660 933 760 977
rect 1008 940 1108 984
rect 1212 940 1312 984
rect 1416 940 1516 984
rect 146 512 246 573
rect 146 466 187 512
rect 233 466 246 512
rect 350 532 450 573
rect 350 486 366 532
rect 412 513 450 532
rect 660 529 760 573
rect 412 486 614 513
rect 350 473 614 486
rect 146 377 246 466
rect 126 333 246 377
rect 350 412 470 425
rect 350 366 363 412
rect 409 366 470 412
rect 350 333 470 366
rect 574 377 614 473
rect 673 483 686 529
rect 732 483 760 529
rect 673 470 760 483
rect 1008 503 1108 580
rect 1008 457 1036 503
rect 1082 457 1108 503
rect 1212 547 1312 580
rect 1212 501 1225 547
rect 1271 520 1312 547
rect 1416 520 1516 580
rect 1271 501 1516 520
rect 1212 480 1516 501
rect 574 333 694 377
rect 1008 376 1108 457
rect 988 332 1108 376
rect 1212 411 1556 432
rect 1212 365 1225 411
rect 1271 392 1556 411
rect 1271 365 1332 392
rect 1212 332 1332 365
rect 1436 332 1556 392
rect 126 25 246 69
rect 350 25 470 69
rect 574 25 694 69
rect 988 24 1108 68
rect 1212 24 1332 68
rect 1436 24 1556 68
<< polycontact >>
rect 187 466 233 512
rect 366 486 412 532
rect 363 366 409 412
rect 686 483 732 529
rect 1036 457 1082 503
rect 1225 501 1271 547
rect 1225 365 1271 411
<< metal1 >>
rect 0 927 1680 1098
rect 0 920 1137 927
rect 0 918 275 920
rect 321 918 1137 920
rect 275 769 321 780
rect 1183 918 1545 927
rect 1137 776 1183 787
rect 1591 918 1680 927
rect 1545 776 1591 787
rect 51 726 117 737
rect 51 586 71 726
rect 51 412 117 586
rect 585 726 978 737
rect 631 701 978 726
rect 1341 733 1426 744
rect 631 691 1271 701
rect 933 655 1271 691
rect 585 575 631 586
rect 789 632 835 643
rect 176 532 418 543
rect 176 512 366 532
rect 176 466 187 512
rect 233 486 366 512
rect 412 486 418 532
rect 233 466 418 486
rect 464 483 686 529
rect 732 483 743 529
rect 464 412 510 483
rect 789 437 835 586
rect 51 366 363 412
rect 409 366 510 412
rect 631 391 835 437
rect 933 639 979 655
rect 51 320 97 366
rect 631 298 677 391
rect 933 331 979 593
rect 1225 547 1271 655
rect 1025 503 1093 542
rect 1025 457 1036 503
rect 1082 457 1093 503
rect 1225 490 1271 501
rect 1387 593 1426 733
rect 499 287 677 298
rect 51 169 97 180
rect 275 222 321 233
rect 0 82 275 90
rect 545 217 677 287
rect 723 320 979 331
rect 769 274 979 320
rect 723 263 979 274
rect 1025 365 1225 411
rect 1271 365 1282 411
rect 1025 217 1071 365
rect 1341 319 1426 593
rect 545 206 1071 217
rect 545 160 913 206
rect 959 160 1071 206
rect 545 147 1071 160
rect 499 136 1071 147
rect 1137 221 1183 232
rect 321 82 1137 90
rect 0 81 1137 82
rect 1341 179 1361 319
rect 1407 179 1426 319
rect 1341 168 1426 179
rect 1585 221 1631 232
rect 1183 81 1585 90
rect 1631 81 1680 90
rect 0 -90 1680 81
<< labels >>
flabel metal1 s 176 466 418 543 0 FreeSans 200 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1025 457 1093 542 0 FreeSans 200 0 0 0 I
port 2 nsew default input
flabel metal1 s 0 918 1680 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 275 232 321 233 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 1341 168 1426 744 0 FreeSans 200 0 0 0 Z
port 3 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 1545 776 1591 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1137 776 1183 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 275 776 321 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 275 769 321 776 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1585 90 1631 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1137 90 1183 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 275 90 321 232 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1680 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1680 1008
string GDS_END 1309858
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1304702
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
