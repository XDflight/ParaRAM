magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -205 231 205 236
rect -205 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 205 231
rect -205 169 205 203
rect -205 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 205 169
rect -205 107 205 141
rect -205 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 205 107
rect -205 45 205 79
rect -205 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 205 45
rect -205 -17 205 17
rect -205 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 205 -17
rect -205 -79 205 -45
rect -205 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 205 -79
rect -205 -141 205 -107
rect -205 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 205 -141
rect -205 -203 205 -169
rect -205 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 205 -203
rect -205 -236 205 -231
<< via2 >>
rect -200 203 -172 231
rect -138 203 -110 231
rect -76 203 -48 231
rect -14 203 14 231
rect 48 203 76 231
rect 110 203 138 231
rect 172 203 200 231
rect -200 141 -172 169
rect -138 141 -110 169
rect -76 141 -48 169
rect -14 141 14 169
rect 48 141 76 169
rect 110 141 138 169
rect 172 141 200 169
rect -200 79 -172 107
rect -138 79 -110 107
rect -76 79 -48 107
rect -14 79 14 107
rect 48 79 76 107
rect 110 79 138 107
rect 172 79 200 107
rect -200 17 -172 45
rect -138 17 -110 45
rect -76 17 -48 45
rect -14 17 14 45
rect 48 17 76 45
rect 110 17 138 45
rect 172 17 200 45
rect -200 -45 -172 -17
rect -138 -45 -110 -17
rect -76 -45 -48 -17
rect -14 -45 14 -17
rect 48 -45 76 -17
rect 110 -45 138 -17
rect 172 -45 200 -17
rect -200 -107 -172 -79
rect -138 -107 -110 -79
rect -76 -107 -48 -79
rect -14 -107 14 -79
rect 48 -107 76 -79
rect 110 -107 138 -79
rect 172 -107 200 -79
rect -200 -169 -172 -141
rect -138 -169 -110 -141
rect -76 -169 -48 -141
rect -14 -169 14 -141
rect 48 -169 76 -141
rect 110 -169 138 -141
rect 172 -169 200 -141
rect -200 -231 -172 -203
rect -138 -231 -110 -203
rect -76 -231 -48 -203
rect -14 -231 14 -203
rect 48 -231 76 -203
rect 110 -231 138 -203
rect 172 -231 200 -203
<< metal3 >>
rect -205 231 205 236
rect -205 203 -200 231
rect -172 203 -138 231
rect -110 203 -76 231
rect -48 203 -14 231
rect 14 203 48 231
rect 76 203 110 231
rect 138 203 172 231
rect 200 203 205 231
rect -205 169 205 203
rect -205 141 -200 169
rect -172 141 -138 169
rect -110 141 -76 169
rect -48 141 -14 169
rect 14 141 48 169
rect 76 141 110 169
rect 138 141 172 169
rect 200 141 205 169
rect -205 107 205 141
rect -205 79 -200 107
rect -172 79 -138 107
rect -110 79 -76 107
rect -48 79 -14 107
rect 14 79 48 107
rect 76 79 110 107
rect 138 79 172 107
rect 200 79 205 107
rect -205 45 205 79
rect -205 17 -200 45
rect -172 17 -138 45
rect -110 17 -76 45
rect -48 17 -14 45
rect 14 17 48 45
rect 76 17 110 45
rect 138 17 172 45
rect 200 17 205 45
rect -205 -17 205 17
rect -205 -45 -200 -17
rect -172 -45 -138 -17
rect -110 -45 -76 -17
rect -48 -45 -14 -17
rect 14 -45 48 -17
rect 76 -45 110 -17
rect 138 -45 172 -17
rect 200 -45 205 -17
rect -205 -79 205 -45
rect -205 -107 -200 -79
rect -172 -107 -138 -79
rect -110 -107 -76 -79
rect -48 -107 -14 -79
rect 14 -107 48 -79
rect 76 -107 110 -79
rect 138 -107 172 -79
rect 200 -107 205 -79
rect -205 -141 205 -107
rect -205 -169 -200 -141
rect -172 -169 -138 -141
rect -110 -169 -76 -141
rect -48 -169 -14 -141
rect 14 -169 48 -141
rect 76 -169 110 -141
rect 138 -169 172 -141
rect 200 -169 205 -141
rect -205 -203 205 -169
rect -205 -231 -200 -203
rect -172 -231 -138 -203
rect -110 -231 -76 -203
rect -48 -231 -14 -203
rect 14 -231 48 -203
rect 76 -231 110 -203
rect 138 -231 172 -203
rect 200 -231 205 -203
rect -205 -236 205 -231
<< properties >>
string GDS_END 1146046
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1142330
<< end >>
