magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 323 29342 342
rect -42 -23 -23 323
rect 29323 -23 29342 323
rect -42 -42 29342 -23
<< psubdiffcont >>
rect -23 -23 29323 323
<< metal1 >>
rect -34 323 29334 334
rect -34 -23 -23 323
rect 29323 -23 29334 323
rect -34 -34 29334 -23
<< properties >>
string GDS_END 1242544
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1167084
<< end >>
