magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1430 1094
<< pwell >>
rect -86 -86 1430 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 806 573 906 939
rect 1020 573 1120 939
<< mvndiff >>
rect 36 305 124 333
rect 36 165 49 305
rect 95 165 124 305
rect 36 69 124 165
rect 244 305 348 333
rect 244 165 273 305
rect 319 165 348 305
rect 244 69 348 165
rect 468 305 572 333
rect 468 165 497 305
rect 543 165 572 305
rect 468 69 572 165
rect 692 305 796 333
rect 692 165 721 305
rect 767 165 796 305
rect 692 69 796 165
rect 916 285 1020 333
rect 916 239 945 285
rect 991 239 1020 285
rect 916 69 1020 239
rect 1140 305 1228 333
rect 1140 165 1169 305
rect 1215 165 1228 305
rect 1140 69 1228 165
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 573 582 939
rect 682 861 806 939
rect 682 721 731 861
rect 777 721 806 861
rect 682 573 806 721
rect 906 573 1020 939
rect 1120 861 1208 939
rect 1120 721 1149 861
rect 1195 721 1208 861
rect 1120 573 1208 721
<< mvndiffc >>
rect 49 165 95 305
rect 273 165 319 305
rect 497 165 543 305
rect 721 165 767 305
rect 945 239 991 285
rect 1169 165 1215 305
<< mvpdiffc >>
rect 69 721 115 861
rect 731 721 777 861
rect 1149 721 1195 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 806 939 906 983
rect 1020 939 1120 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 377 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 377 458 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 377 682 454
rect 806 500 906 573
rect 806 454 819 500
rect 865 454 906 500
rect 806 377 906 454
rect 1020 500 1120 573
rect 1020 454 1038 500
rect 1084 454 1120 500
rect 1020 377 1120 454
rect 124 333 244 377
rect 348 333 468 377
rect 572 333 692 377
rect 796 333 916 377
rect 1020 333 1140 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 595 454 641 500
rect 819 454 865 500
rect 1038 454 1084 500
<< metal1 >>
rect 0 918 1344 1098
rect 69 861 115 918
rect 69 710 115 721
rect 731 861 777 872
rect 731 603 777 721
rect 1149 861 1195 918
rect 1149 710 1195 721
rect 731 557 991 603
rect 142 500 203 542
rect 142 454 157 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 584 500 652 542
rect 584 454 595 500
rect 641 454 652 500
rect 814 500 866 511
rect 814 454 819 500
rect 865 454 866 500
rect 142 443 203 454
rect 273 362 767 408
rect 49 305 95 316
rect 49 90 95 165
rect 273 305 319 362
rect 273 154 319 165
rect 497 305 543 316
rect 497 90 543 165
rect 721 305 767 362
rect 814 354 866 454
rect 926 285 991 557
rect 1038 500 1090 511
rect 1084 454 1090 500
rect 1038 354 1090 454
rect 926 239 945 285
rect 926 228 991 239
rect 1169 305 1215 316
rect 767 165 1169 182
rect 721 136 1215 165
rect 0 -90 1344 90
<< labels >>
flabel metal1 s 584 454 652 542 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 142 443 203 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 814 354 866 511 0 FreeSans 200 0 0 0 B1
port 4 nsew default input
flabel metal1 s 1038 354 1090 511 0 FreeSans 200 0 0 0 B2
port 5 nsew default input
flabel metal1 s 0 918 1344 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 497 90 543 316 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 731 603 777 872 0 FreeSans 200 0 0 0 ZN
port 6 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 731 557 991 603 1 ZN
port 6 nsew default output
rlabel metal1 s 926 228 991 557 1 ZN
port 6 nsew default output
rlabel metal1 s 1149 710 1195 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 49 90 95 316 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 1344 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1344 1008
string GDS_END 162176
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 158114
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
