magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 776 1028
<< mvpmos >>
rect 0 0 120 908
rect 224 0 344 908
rect 448 0 568 908
<< mvpdiff >>
rect -88 895 0 908
rect -88 849 -75 895
rect -29 849 0 895
rect -88 791 0 849
rect -88 745 -75 791
rect -29 745 0 791
rect -88 687 0 745
rect -88 641 -75 687
rect -29 641 0 687
rect -88 583 0 641
rect -88 537 -75 583
rect -29 537 0 583
rect -88 479 0 537
rect -88 433 -75 479
rect -29 433 0 479
rect -88 374 0 433
rect -88 328 -75 374
rect -29 328 0 374
rect -88 269 0 328
rect -88 223 -75 269
rect -29 223 0 269
rect -88 164 0 223
rect -88 118 -75 164
rect -29 118 0 164
rect -88 59 0 118
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 895 224 908
rect 120 849 149 895
rect 195 849 224 895
rect 120 791 224 849
rect 120 745 149 791
rect 195 745 224 791
rect 120 687 224 745
rect 120 641 149 687
rect 195 641 224 687
rect 120 583 224 641
rect 120 537 149 583
rect 195 537 224 583
rect 120 479 224 537
rect 120 433 149 479
rect 195 433 224 479
rect 120 374 224 433
rect 120 328 149 374
rect 195 328 224 374
rect 120 269 224 328
rect 120 223 149 269
rect 195 223 224 269
rect 120 164 224 223
rect 120 118 149 164
rect 195 118 224 164
rect 120 59 224 118
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 895 448 908
rect 344 849 373 895
rect 419 849 448 895
rect 344 791 448 849
rect 344 745 373 791
rect 419 745 448 791
rect 344 687 448 745
rect 344 641 373 687
rect 419 641 448 687
rect 344 583 448 641
rect 344 537 373 583
rect 419 537 448 583
rect 344 479 448 537
rect 344 433 373 479
rect 419 433 448 479
rect 344 374 448 433
rect 344 328 373 374
rect 419 328 448 374
rect 344 269 448 328
rect 344 223 373 269
rect 419 223 448 269
rect 344 164 448 223
rect 344 118 373 164
rect 419 118 448 164
rect 344 59 448 118
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 895 656 908
rect 568 849 597 895
rect 643 849 656 895
rect 568 791 656 849
rect 568 745 597 791
rect 643 745 656 791
rect 568 687 656 745
rect 568 641 597 687
rect 643 641 656 687
rect 568 583 656 641
rect 568 537 597 583
rect 643 537 656 583
rect 568 479 656 537
rect 568 433 597 479
rect 643 433 656 479
rect 568 374 656 433
rect 568 328 597 374
rect 643 328 656 374
rect 568 269 656 328
rect 568 223 597 269
rect 643 223 656 269
rect 568 164 656 223
rect 568 118 597 164
rect 643 118 656 164
rect 568 59 656 118
rect 568 13 597 59
rect 643 13 656 59
rect 568 0 656 13
<< mvpdiffc >>
rect -75 849 -29 895
rect -75 745 -29 791
rect -75 641 -29 687
rect -75 537 -29 583
rect -75 433 -29 479
rect -75 328 -29 374
rect -75 223 -29 269
rect -75 118 -29 164
rect -75 13 -29 59
rect 149 849 195 895
rect 149 745 195 791
rect 149 641 195 687
rect 149 537 195 583
rect 149 433 195 479
rect 149 328 195 374
rect 149 223 195 269
rect 149 118 195 164
rect 149 13 195 59
rect 373 849 419 895
rect 373 745 419 791
rect 373 641 419 687
rect 373 537 419 583
rect 373 433 419 479
rect 373 328 419 374
rect 373 223 419 269
rect 373 118 419 164
rect 373 13 419 59
rect 597 849 643 895
rect 597 745 643 791
rect 597 641 643 687
rect 597 537 643 583
rect 597 433 643 479
rect 597 328 643 374
rect 597 223 643 269
rect 597 118 643 164
rect 597 13 643 59
<< polysilicon >>
rect 0 908 120 952
rect 224 908 344 952
rect 448 908 568 952
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
<< metal1 >>
rect -75 895 -29 908
rect -75 791 -29 849
rect -75 687 -29 745
rect -75 583 -29 641
rect -75 479 -29 537
rect -75 374 -29 433
rect -75 269 -29 328
rect -75 164 -29 223
rect -75 59 -29 118
rect -75 0 -29 13
rect 149 895 195 908
rect 149 791 195 849
rect 149 687 195 745
rect 149 583 195 641
rect 149 479 195 537
rect 149 374 195 433
rect 149 269 195 328
rect 149 164 195 223
rect 149 59 195 118
rect 149 0 195 13
rect 373 895 419 908
rect 373 791 419 849
rect 373 687 419 745
rect 373 583 419 641
rect 373 479 419 537
rect 373 374 419 433
rect 373 269 419 328
rect 373 164 419 223
rect 373 59 419 118
rect 373 0 419 13
rect 597 895 643 908
rect 597 791 643 849
rect 597 687 643 745
rect 597 583 643 641
rect 597 479 643 537
rect 597 374 643 433
rect 597 269 643 328
rect 597 164 643 223
rect 597 59 643 118
rect 597 0 643 13
<< labels >>
flabel metal1 s -52 454 -52 454 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 454 620 454 0 FreeSans 400 0 0 0 D
flabel metal1 s 172 454 172 454 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 454 396 454 0 FreeSans 400 0 0 0 S
<< properties >>
string GDS_END 116798
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 112770
<< end >>
