magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 462 4342 1094
rect -86 453 86 462
rect 3842 454 4342 462
rect 4170 453 4342 454
<< pwell >>
rect 1854 453 3542 462
rect -86 -86 4342 453
<< mvnmos >>
rect 124 156 244 272
rect 348 156 468 272
rect 516 156 636 272
rect 740 156 860 272
rect 908 156 1028 272
rect 1308 156 1428 314
rect 1620 156 1740 314
rect 1988 226 2108 342
rect 2212 226 2332 342
rect 2380 226 2500 342
rect 2680 226 2800 342
rect 2904 226 3024 342
rect 3128 226 3248 342
rect 3296 226 3416 342
rect 3596 183 3716 333
rect 3964 69 4084 333
<< mvpmos >>
rect 134 652 234 852
rect 345 652 445 852
rect 496 652 596 852
rect 700 652 800 852
rect 888 652 988 852
rect 1318 582 1418 858
rect 1612 582 1712 858
rect 1998 652 2098 852
rect 2212 652 2312 852
rect 2390 652 2490 852
rect 2674 652 2774 852
rect 2914 652 3014 852
rect 3128 652 3228 852
rect 3276 652 3376 852
rect 3516 632 3616 852
rect 3974 574 4074 940
<< mvndiff >>
rect 1220 297 1308 314
rect 36 215 124 272
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 272
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 272
rect 636 215 740 272
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 272
rect 1028 156 1148 272
rect 1220 251 1233 297
rect 1279 251 1308 297
rect 1220 156 1308 251
rect 1428 156 1620 314
rect 1740 301 1828 314
rect 1740 255 1769 301
rect 1815 255 1828 301
rect 1740 156 1828 255
rect 1900 285 1988 342
rect 1900 239 1913 285
rect 1959 239 1988 285
rect 1900 226 1988 239
rect 2108 329 2212 342
rect 2108 283 2137 329
rect 2183 283 2212 329
rect 2108 226 2212 283
rect 2332 226 2380 342
rect 2500 226 2680 342
rect 2800 329 2904 342
rect 2800 283 2829 329
rect 2875 283 2904 329
rect 2800 226 2904 283
rect 3024 329 3128 342
rect 3024 283 3053 329
rect 3099 283 3128 329
rect 3024 226 3128 283
rect 3248 226 3296 342
rect 3416 333 3496 342
rect 3416 226 3596 333
rect 1088 115 1148 156
rect 1088 102 1160 115
rect 1088 56 1101 102
rect 1147 56 1160 102
rect 1088 43 1160 56
rect 1488 102 1560 156
rect 1488 56 1501 102
rect 1547 56 1560 102
rect 1488 43 1560 56
rect 2560 114 2620 226
rect 3476 183 3596 226
rect 3716 320 3804 333
rect 3716 274 3745 320
rect 3791 274 3804 320
rect 3716 183 3804 274
rect 3876 309 3964 333
rect 3476 146 3536 183
rect 3464 133 3536 146
rect 3876 169 3889 309
rect 3935 169 3964 309
rect 2560 101 2632 114
rect 2560 55 2573 101
rect 2619 55 2632 101
rect 3464 87 3477 133
rect 3523 87 3536 133
rect 3464 74 3536 87
rect 3876 69 3964 169
rect 4084 309 4172 333
rect 4084 169 4113 309
rect 4159 169 4172 309
rect 4084 69 4172 169
rect 2560 42 2632 55
<< mvpdiff >>
rect 46 839 134 852
rect 46 699 59 839
rect 105 699 134 839
rect 46 652 134 699
rect 234 839 345 852
rect 234 699 263 839
rect 309 699 345 839
rect 234 652 345 699
rect 445 652 496 852
rect 596 839 700 852
rect 596 699 625 839
rect 671 699 700 839
rect 596 652 700 699
rect 800 652 888 852
rect 988 839 1076 852
rect 988 793 1017 839
rect 1063 793 1076 839
rect 988 652 1076 793
rect 1193 644 1318 858
rect 1193 598 1206 644
rect 1252 598 1318 644
rect 1193 582 1318 598
rect 1418 845 1612 858
rect 1418 799 1447 845
rect 1493 799 1612 845
rect 1418 582 1612 799
rect 1712 641 1800 858
rect 1910 758 1998 852
rect 1910 712 1923 758
rect 1969 712 1998 758
rect 1910 652 1998 712
rect 2098 839 2212 852
rect 2098 699 2137 839
rect 2183 699 2212 839
rect 2098 652 2212 699
rect 2312 652 2390 852
rect 2490 839 2674 852
rect 2490 699 2519 839
rect 2565 699 2674 839
rect 2490 652 2674 699
rect 2774 839 2914 852
rect 2774 699 2803 839
rect 2849 699 2914 839
rect 2774 652 2914 699
rect 3014 839 3128 852
rect 3014 699 3053 839
rect 3099 699 3128 839
rect 3014 652 3128 699
rect 3228 652 3276 852
rect 3376 776 3516 852
rect 3376 730 3405 776
rect 3451 730 3516 776
rect 3376 652 3516 730
rect 1712 595 1741 641
rect 1787 595 1800 641
rect 1712 582 1800 595
rect 3436 632 3516 652
rect 3616 839 3704 852
rect 3616 699 3645 839
rect 3691 699 3704 839
rect 3616 632 3704 699
rect 3886 727 3974 940
rect 3886 587 3899 727
rect 3945 587 3974 727
rect 3886 574 3974 587
rect 4074 927 4162 940
rect 4074 787 4103 927
rect 4149 787 4162 927
rect 4074 574 4162 787
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1233 251 1279 297
rect 1769 255 1815 301
rect 1913 239 1959 285
rect 2137 283 2183 329
rect 2829 283 2875 329
rect 3053 283 3099 329
rect 1101 56 1147 102
rect 1501 56 1547 102
rect 3745 274 3791 320
rect 3889 169 3935 309
rect 2573 55 2619 101
rect 3477 87 3523 133
rect 4113 169 4159 309
<< mvpdiffc >>
rect 59 699 105 839
rect 263 699 309 839
rect 625 699 671 839
rect 1017 793 1063 839
rect 1206 598 1252 644
rect 1447 799 1493 845
rect 1923 712 1969 758
rect 2137 699 2183 839
rect 2519 699 2565 839
rect 2803 699 2849 839
rect 3053 699 3099 839
rect 3405 730 3451 776
rect 1741 595 1787 641
rect 3645 699 3691 839
rect 3899 587 3945 727
rect 4103 787 4149 927
<< polysilicon >>
rect 134 944 800 984
rect 134 852 234 944
rect 345 852 445 896
rect 496 852 596 896
rect 700 852 800 944
rect 1612 944 3014 984
rect 888 852 988 896
rect 1318 858 1418 902
rect 1612 858 1712 944
rect 134 506 234 652
rect 124 493 234 506
rect 124 447 137 493
rect 183 447 234 493
rect 124 316 234 447
rect 345 493 445 652
rect 345 447 358 493
rect 404 447 445 493
rect 345 439 445 447
rect 348 316 445 439
rect 496 493 596 652
rect 700 608 800 652
rect 888 608 988 652
rect 496 447 509 493
rect 555 447 596 493
rect 496 436 596 447
rect 908 493 988 608
rect 1998 852 2098 896
rect 2212 852 2312 944
rect 2390 852 2490 896
rect 2674 852 2774 896
rect 2914 852 3014 944
rect 3974 940 4074 984
rect 3128 852 3228 896
rect 3276 852 3376 896
rect 3516 852 3616 896
rect 1318 506 1418 582
rect 908 447 926 493
rect 972 447 988 493
rect 496 364 860 436
rect 124 272 244 316
rect 348 272 468 316
rect 516 272 636 316
rect 740 272 860 364
rect 908 316 988 447
rect 1308 493 1418 506
rect 1308 447 1321 493
rect 1367 447 1418 493
rect 1308 358 1418 447
rect 1612 493 1712 582
rect 1612 447 1625 493
rect 1671 447 1712 493
rect 1612 435 1712 447
rect 1620 358 1712 435
rect 1998 506 2098 652
rect 2212 608 2312 652
rect 2390 506 2490 652
rect 1998 493 2332 506
rect 1998 447 2011 493
rect 2057 447 2332 493
rect 1998 434 2332 447
rect 908 272 1028 316
rect 1308 314 1428 358
rect 1620 314 1740 358
rect 1988 342 2108 386
rect 2212 342 2332 434
rect 2390 493 2500 506
rect 2390 447 2441 493
rect 2487 447 2500 493
rect 2390 386 2500 447
rect 2674 493 2774 652
rect 2674 447 2687 493
rect 2733 447 2774 493
rect 2674 436 2774 447
rect 2380 342 2500 386
rect 2680 386 2774 436
rect 2914 474 3014 652
rect 3128 581 3228 652
rect 3276 608 3376 652
rect 3128 535 3156 581
rect 3202 535 3228 581
rect 3128 522 3228 535
rect 3296 506 3376 608
rect 3296 493 3416 506
rect 2914 434 3248 474
rect 2680 342 2800 386
rect 2904 342 3024 386
rect 3128 342 3248 434
rect 3296 447 3337 493
rect 3383 447 3416 493
rect 3296 342 3416 447
rect 3516 493 3616 632
rect 3974 506 4074 574
rect 3516 447 3529 493
rect 3575 476 3616 493
rect 3732 493 4074 506
rect 3575 447 3656 476
rect 3516 434 3656 447
rect 3732 447 3745 493
rect 3791 447 4074 493
rect 3732 434 4074 447
rect 3596 377 3656 434
rect 3964 377 4074 434
rect 3596 333 3716 377
rect 3964 333 4084 377
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 124 24 636 64
rect 1308 112 1428 156
rect 1620 96 1740 156
rect 1988 96 2108 226
rect 2212 193 2332 226
rect 2212 147 2273 193
rect 2319 147 2332 193
rect 2380 182 2500 226
rect 2212 134 2332 147
rect 1620 24 2108 96
rect 2680 182 2800 226
rect 2904 193 3024 226
rect 2904 147 2917 193
rect 2963 147 3024 193
rect 3128 182 3248 226
rect 3296 182 3416 226
rect 2904 134 3024 147
rect 3596 139 3716 183
rect 3964 25 4084 69
<< polycontact >>
rect 137 447 183 493
rect 358 447 404 493
rect 509 447 555 493
rect 926 447 972 493
rect 1321 447 1367 493
rect 1625 447 1671 493
rect 2011 447 2057 493
rect 2441 447 2487 493
rect 2687 447 2733 493
rect 3156 535 3202 581
rect 3337 447 3383 493
rect 3529 447 3575 493
rect 3745 447 3791 493
rect 2273 147 2319 193
rect 2917 147 2963 193
<< metal1 >>
rect 0 927 4256 1098
rect 0 918 4103 927
rect 59 839 105 850
rect 59 642 105 699
rect 263 839 309 918
rect 263 688 309 699
rect 625 839 671 850
rect 1006 839 1074 918
rect 1006 793 1017 839
rect 1063 793 1074 839
rect 1436 845 1504 918
rect 1436 799 1447 845
rect 1493 799 1504 845
rect 2137 839 2183 850
rect 1923 758 1969 769
rect 671 712 1923 747
rect 671 701 1969 712
rect 625 688 671 699
rect 1206 644 1671 655
rect 59 596 555 642
rect 30 493 183 542
rect 30 447 137 493
rect 30 436 183 447
rect 254 493 404 542
rect 254 447 358 493
rect 254 436 404 447
rect 509 493 555 596
rect 1252 609 1671 644
rect 1206 587 1252 598
rect 30 354 82 436
rect 254 354 306 436
rect 509 307 555 447
rect 49 261 555 307
rect 926 493 978 504
rect 972 447 978 493
rect 49 215 95 261
rect 926 242 978 447
rect 1262 493 1367 542
rect 1262 447 1321 493
rect 1262 354 1367 447
rect 1625 493 1671 609
rect 1625 308 1671 447
rect 1233 297 1671 308
rect 1279 251 1671 297
rect 1233 240 1671 251
rect 1741 641 1787 652
rect 1741 504 1787 595
rect 1741 493 2057 504
rect 1741 447 2011 493
rect 1741 436 2057 447
rect 1741 301 1815 436
rect 1741 255 1769 301
rect 2137 390 2183 699
rect 2519 839 2565 918
rect 2519 688 2565 699
rect 2803 839 2875 850
rect 2849 699 2875 839
rect 2803 596 2875 699
rect 2441 550 2875 596
rect 2441 493 2487 550
rect 2441 436 2487 447
rect 2687 493 2733 504
rect 2687 390 2733 447
rect 2137 344 2733 390
rect 2137 329 2183 344
rect 1741 244 1815 255
rect 1913 285 1959 296
rect 2137 272 2183 283
rect 2829 329 2875 550
rect 2829 272 2875 283
rect 3053 839 3099 850
rect 3405 776 3451 918
rect 3405 719 3451 730
rect 3645 839 3691 850
rect 3053 673 3099 699
rect 4149 918 4256 927
rect 4103 776 4149 787
rect 3053 627 3586 673
rect 3053 329 3099 627
rect 3053 272 3099 283
rect 3145 535 3156 581
rect 3202 535 3213 581
rect 665 215 711 226
rect 49 158 95 169
rect 262 169 273 215
rect 319 169 330 215
rect 262 90 330 169
rect 1913 194 1959 239
rect 3145 204 3213 535
rect 3518 493 3586 627
rect 3326 447 3337 493
rect 3383 447 3394 493
rect 3518 447 3529 493
rect 3575 447 3586 493
rect 3645 504 3691 699
rect 3899 727 3945 738
rect 3899 542 3945 587
rect 3645 493 3791 504
rect 3645 458 3745 493
rect 3326 309 3394 447
rect 3745 320 3791 447
rect 3326 274 3745 309
rect 3326 263 3791 274
rect 3838 309 3945 542
rect 3838 242 3889 309
rect 711 169 1959 194
rect 665 148 1959 169
rect 2273 193 3213 204
rect 2319 147 2917 193
rect 2963 147 3213 193
rect 3935 169 3945 309
rect 3889 158 3945 169
rect 4113 309 4159 320
rect 2273 136 2319 147
rect 3477 133 3523 144
rect 1090 90 1101 102
rect 0 56 1101 90
rect 1147 90 1158 102
rect 1490 90 1501 102
rect 1147 56 1501 90
rect 1547 90 1558 102
rect 2562 90 2573 101
rect 1547 56 2573 90
rect 0 55 2573 56
rect 2619 90 2630 101
rect 2619 87 3477 90
rect 4113 90 4159 169
rect 3523 87 4256 90
rect 2619 55 4256 87
rect 0 -90 4256 55
<< labels >>
flabel metal1 s 1262 354 1367 542 0 FreeSans 200 0 0 0 CLK
port 4 nsew clock input
flabel metal1 s 926 242 978 504 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 3899 542 3945 738 0 FreeSans 200 0 0 0 Q
port 5 nsew default output
flabel metal1 s 30 436 183 542 0 FreeSans 200 0 0 0 SE
port 2 nsew default input
flabel metal1 s 254 436 404 542 0 FreeSans 200 0 0 0 SI
port 3 nsew default input
flabel metal1 s 0 918 4256 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 4113 215 4159 320 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 30 354 82 436 1 SE
port 2 nsew default input
rlabel metal1 s 254 354 306 436 1 SI
port 3 nsew default input
rlabel metal1 s 3838 242 3945 542 1 Q
port 5 nsew default output
rlabel metal1 s 3889 158 3945 242 1 Q
port 5 nsew default output
rlabel metal1 s 4103 799 4149 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3405 799 3451 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2519 799 2565 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1436 799 1504 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1006 799 1074 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 263 799 309 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4103 793 4149 799 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3405 793 3451 799 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2519 793 2565 799 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1006 793 1074 799 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 263 793 309 799 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4103 776 4149 793 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3405 776 3451 793 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2519 776 2565 793 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 263 776 309 793 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3405 719 3451 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2519 719 2565 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 263 719 309 776 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2519 688 2565 719 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 263 688 309 719 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4113 144 4159 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 144 330 215 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 102 4159 144 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3477 102 3523 144 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 102 330 144 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 101 4159 102 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3477 101 3523 102 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1490 101 1558 102 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1090 101 1158 102 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 101 330 102 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4113 90 4159 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3477 90 3523 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2562 90 2630 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1490 90 1558 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1090 90 1158 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 101 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4256 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 1008
string GDS_END 305490
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 296208
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
