magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -2294 82 -2133 83
rect 1976 82 2294 83
rect -2294 23 2294 82
rect -2294 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 2294 23
rect -2294 -83 2294 -23
<< psubdiffcont >>
rect -1920 -23 -1874 23
rect -1762 -23 -1716 23
rect -1604 -23 -1558 23
rect -1446 -23 -1400 23
rect -1288 -23 -1242 23
rect -1130 -23 -1084 23
rect -972 -23 -926 23
rect -814 -23 -768 23
rect -656 -23 -610 23
rect -497 -23 -451 23
rect -339 -23 -293 23
rect -181 -23 -135 23
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect 1242 -23 1288 23
rect 1400 -23 1446 23
rect 1558 -23 1604 23
rect 1716 -23 1762 23
rect 1874 -23 1920 23
<< metal1 >>
rect -2285 73 -1788 74
rect -705 73 -589 74
rect 191 73 307 74
rect 580 73 696 74
rect 1475 73 2285 74
rect -2285 23 2285 73
rect -2285 -23 -1920 23
rect -1874 -23 -1762 23
rect -1716 -23 -1604 23
rect -1558 -23 -1446 23
rect -1400 -23 -1288 23
rect -1242 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1874 23
rect 1920 -23 2285 23
rect -2285 -74 2285 -23
<< properties >>
string GDS_END 825930
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 823974
<< end >>
