magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 3808 844
rect 49 536 95 724
rect 273 600 319 678
rect 477 646 523 724
rect 701 600 747 678
rect 925 646 971 724
rect 1149 600 1195 678
rect 1373 646 1419 724
rect 1616 600 1662 678
rect 1821 646 1867 724
rect 2045 600 2091 678
rect 2269 646 2315 724
rect 2493 600 2539 678
rect 2717 646 2763 724
rect 2941 600 2987 678
rect 3165 646 3211 724
rect 3389 600 3435 678
rect 273 484 3435 600
rect 3613 536 3659 724
rect 124 353 1702 438
rect 1758 289 1938 484
rect 2003 353 3584 438
rect 49 60 95 203
rect 273 173 3455 289
rect 273 135 325 173
rect 721 135 767 173
rect 1169 135 1215 173
rect 1617 135 1663 173
rect 2065 135 2111 173
rect 2513 135 2559 173
rect 2961 135 3007 173
rect 3409 135 3455 173
rect 486 60 554 127
rect 934 60 1002 127
rect 1382 60 1450 127
rect 1830 60 1898 127
rect 2278 60 2346 127
rect 2726 60 2794 127
rect 3174 60 3242 127
rect 3633 60 3679 203
rect 0 -60 3808 60
<< labels >>
rlabel metal1 s 124 353 1702 438 6 I
port 1 nsew default input
rlabel metal1 s 2003 353 3584 438 6 I
port 1 nsew default input
rlabel metal1 s 3389 600 3435 678 6 ZN
port 2 nsew default output
rlabel metal1 s 2941 600 2987 678 6 ZN
port 2 nsew default output
rlabel metal1 s 2493 600 2539 678 6 ZN
port 2 nsew default output
rlabel metal1 s 2045 600 2091 678 6 ZN
port 2 nsew default output
rlabel metal1 s 1616 600 1662 678 6 ZN
port 2 nsew default output
rlabel metal1 s 1149 600 1195 678 6 ZN
port 2 nsew default output
rlabel metal1 s 701 600 747 678 6 ZN
port 2 nsew default output
rlabel metal1 s 273 600 319 678 6 ZN
port 2 nsew default output
rlabel metal1 s 273 484 3435 600 6 ZN
port 2 nsew default output
rlabel metal1 s 1758 289 1938 484 6 ZN
port 2 nsew default output
rlabel metal1 s 273 173 3455 289 6 ZN
port 2 nsew default output
rlabel metal1 s 3409 135 3455 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2961 135 3007 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2513 135 2559 173 6 ZN
port 2 nsew default output
rlabel metal1 s 2065 135 2111 173 6 ZN
port 2 nsew default output
rlabel metal1 s 1617 135 1663 173 6 ZN
port 2 nsew default output
rlabel metal1 s 1169 135 1215 173 6 ZN
port 2 nsew default output
rlabel metal1 s 721 135 767 173 6 ZN
port 2 nsew default output
rlabel metal1 s 273 135 325 173 6 ZN
port 2 nsew default output
rlabel metal1 s 0 724 3808 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 646 3659 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 646 3211 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 646 2763 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 646 2315 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 646 1867 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 646 1419 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 646 971 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 646 523 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 646 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 536 3659 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 536 95 646 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3633 127 3679 203 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 127 95 203 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3633 60 3679 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 127 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3808 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 496908
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 488312
<< end >>
