magic
tech gf180mcuC
magscale 1 10
timestamp 1667403444
<< checkpaint >>
rect -2000 -2000 2001 2001
<< end >>
