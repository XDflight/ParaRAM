magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 604
<< mvndiff >>
rect -88 591 0 604
rect -88 545 -75 591
rect -29 545 0 591
rect -88 485 0 545
rect -88 439 -75 485
rect -29 439 0 485
rect -88 379 0 439
rect -88 333 -75 379
rect -29 333 0 379
rect -88 273 0 333
rect -88 227 -75 273
rect -29 227 0 273
rect -88 166 0 227
rect -88 120 -75 166
rect -29 120 0 166
rect -88 59 0 120
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 591 208 604
rect 120 545 149 591
rect 195 545 208 591
rect 120 485 208 545
rect 120 439 149 485
rect 195 439 208 485
rect 120 379 208 439
rect 120 333 149 379
rect 195 333 208 379
rect 120 273 208 333
rect 120 227 149 273
rect 195 227 208 273
rect 120 166 208 227
rect 120 120 149 166
rect 195 120 208 166
rect 120 59 208 120
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 545 -29 591
rect -75 439 -29 485
rect -75 333 -29 379
rect -75 227 -29 273
rect -75 120 -29 166
rect -75 13 -29 59
rect 149 545 195 591
rect 149 439 195 485
rect 149 333 195 379
rect 149 227 195 273
rect 149 120 195 166
rect 149 13 195 59
<< polysilicon >>
rect 0 604 120 648
rect 0 -44 120 0
<< metal1 >>
rect -75 591 -29 604
rect -75 485 -29 545
rect -75 379 -29 439
rect -75 273 -29 333
rect -75 166 -29 227
rect -75 59 -29 120
rect -75 0 -29 13
rect 149 591 195 604
rect 149 485 195 545
rect 149 379 195 439
rect 149 273 195 333
rect 149 166 195 227
rect 149 59 195 120
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 302 -52 302 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 302 172 302 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 591784
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 590120
<< end >>
