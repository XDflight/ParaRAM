magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -170 14063 170 14104
rect -170 14011 -132 14063
rect -80 14011 80 14063
rect 132 14011 170 14063
rect -170 13846 170 14011
rect -170 13794 -132 13846
rect -80 13794 80 13846
rect 132 13794 170 13846
rect -170 13628 170 13794
rect -170 13576 -132 13628
rect -80 13576 80 13628
rect 132 13576 170 13628
rect -170 13410 170 13576
rect -170 13358 -132 13410
rect -80 13358 80 13410
rect 132 13358 170 13410
rect -170 13193 170 13358
rect -170 13141 -132 13193
rect -80 13141 80 13193
rect 132 13141 170 13193
rect -170 12975 170 13141
rect -170 12923 -132 12975
rect -80 12923 80 12975
rect 132 12923 170 12975
rect -170 12758 170 12923
rect -170 12706 -132 12758
rect -80 12706 80 12758
rect 132 12706 170 12758
rect -170 12540 170 12706
rect -170 12488 -132 12540
rect -80 12488 80 12540
rect 132 12488 170 12540
rect -170 12322 170 12488
rect -170 12270 -132 12322
rect -80 12270 80 12322
rect 132 12270 170 12322
rect -170 12105 170 12270
rect -170 12053 -132 12105
rect -80 12053 80 12105
rect 132 12053 170 12105
rect -170 11887 170 12053
rect -170 11835 -132 11887
rect -80 11835 80 11887
rect 132 11835 170 11887
rect -170 11669 170 11835
rect -170 11617 -132 11669
rect -80 11617 80 11669
rect 132 11617 170 11669
rect -170 11452 170 11617
rect -170 11400 -132 11452
rect -80 11400 80 11452
rect 132 11400 170 11452
rect -170 11234 170 11400
rect -170 11182 -132 11234
rect -80 11182 80 11234
rect 132 11182 170 11234
rect -170 11017 170 11182
rect -170 10965 -132 11017
rect -80 10965 80 11017
rect 132 10965 170 11017
rect -170 10799 170 10965
rect -170 10747 -132 10799
rect -80 10747 80 10799
rect 132 10747 170 10799
rect -170 10581 170 10747
rect -170 10529 -132 10581
rect -80 10529 80 10581
rect 132 10529 170 10581
rect -170 10364 170 10529
rect -170 10312 -132 10364
rect -80 10312 80 10364
rect 132 10312 170 10364
rect -170 10146 170 10312
rect -170 10094 -132 10146
rect -80 10094 80 10146
rect 132 10094 170 10146
rect -170 9928 170 10094
rect -170 9876 -132 9928
rect -80 9876 80 9928
rect 132 9876 170 9928
rect -170 9711 170 9876
rect -170 9659 -132 9711
rect -80 9659 80 9711
rect 132 9659 170 9711
rect -170 9493 170 9659
rect -170 9441 -132 9493
rect -80 9441 80 9493
rect 132 9441 170 9493
rect -170 9275 170 9441
rect -170 9223 -132 9275
rect -80 9223 80 9275
rect 132 9223 170 9275
rect -170 9058 170 9223
rect -170 9006 -132 9058
rect -80 9006 80 9058
rect 132 9006 170 9058
rect -170 8840 170 9006
rect -170 8788 -132 8840
rect -80 8788 80 8840
rect 132 8788 170 8840
rect -170 8623 170 8788
rect -170 8571 -132 8623
rect -80 8571 80 8623
rect 132 8571 170 8623
rect -170 8405 170 8571
rect -170 8353 -132 8405
rect -80 8353 80 8405
rect 132 8353 170 8405
rect -170 8187 170 8353
rect -170 8135 -132 8187
rect -80 8135 80 8187
rect 132 8135 170 8187
rect -170 7970 170 8135
rect -170 7918 -132 7970
rect -80 7918 80 7970
rect 132 7918 170 7970
rect -170 7752 170 7918
rect -170 7700 -132 7752
rect -80 7700 80 7752
rect 132 7700 170 7752
rect -170 7534 170 7700
rect -170 7482 -132 7534
rect -80 7482 80 7534
rect 132 7482 170 7534
rect -170 7317 170 7482
rect -170 7265 -132 7317
rect -80 7265 80 7317
rect 132 7265 170 7317
rect -170 7099 170 7265
rect -170 7047 -132 7099
rect -80 7047 80 7099
rect 132 7047 170 7099
rect -170 6881 170 7047
rect -170 6829 -132 6881
rect -80 6829 80 6881
rect 132 6829 170 6881
rect -170 6664 170 6829
rect -170 6612 -132 6664
rect -80 6612 80 6664
rect 132 6612 170 6664
rect -170 6446 170 6612
rect -170 6394 -132 6446
rect -80 6394 80 6446
rect 132 6394 170 6446
rect -170 6229 170 6394
rect -170 6177 -132 6229
rect -80 6177 80 6229
rect 132 6177 170 6229
rect -170 6011 170 6177
rect -170 5959 -132 6011
rect -80 5959 80 6011
rect 132 5959 170 6011
rect -170 5793 170 5959
rect -170 5741 -132 5793
rect -80 5741 80 5793
rect 132 5741 170 5793
rect -170 5576 170 5741
rect -170 5524 -132 5576
rect -80 5524 80 5576
rect 132 5524 170 5576
rect -170 5358 170 5524
rect -170 5306 -132 5358
rect -80 5306 80 5358
rect 132 5306 170 5358
rect -170 5140 170 5306
rect -170 5088 -132 5140
rect -80 5088 80 5140
rect 132 5088 170 5140
rect -170 4923 170 5088
rect -170 4871 -132 4923
rect -80 4871 80 4923
rect 132 4871 170 4923
rect -170 4705 170 4871
rect -170 4653 -132 4705
rect -80 4653 80 4705
rect 132 4653 170 4705
rect -170 4488 170 4653
rect -170 4436 -132 4488
rect -80 4436 80 4488
rect 132 4436 170 4488
rect -170 4270 170 4436
rect -170 4218 -132 4270
rect -80 4218 80 4270
rect 132 4218 170 4270
rect -170 4052 170 4218
rect -170 4000 -132 4052
rect -80 4000 80 4052
rect 132 4000 170 4052
rect -170 3835 170 4000
rect -170 3783 -132 3835
rect -80 3783 80 3835
rect 132 3783 170 3835
rect -170 3617 170 3783
rect -170 3565 -132 3617
rect -80 3565 80 3617
rect 132 3565 170 3617
rect -170 3399 170 3565
rect -170 3347 -132 3399
rect -80 3347 80 3399
rect 132 3347 170 3399
rect -170 3182 170 3347
rect -170 3130 -132 3182
rect -80 3130 80 3182
rect 132 3130 170 3182
rect -170 2964 170 3130
rect -170 2912 -132 2964
rect -80 2912 80 2964
rect 132 2912 170 2964
rect -170 2746 170 2912
rect -170 2694 -132 2746
rect -80 2694 80 2746
rect 132 2694 170 2746
rect -170 2529 170 2694
rect -170 2477 -132 2529
rect -80 2477 80 2529
rect 132 2477 170 2529
rect -170 2311 170 2477
rect -170 2259 -132 2311
rect -80 2259 80 2311
rect 132 2259 170 2311
rect -170 2094 170 2259
rect -170 2042 -132 2094
rect -80 2042 80 2094
rect 132 2042 170 2094
rect -170 1876 170 2042
rect -170 1824 -132 1876
rect -80 1824 80 1876
rect 132 1824 170 1876
rect -170 1658 170 1824
rect -170 1606 -132 1658
rect -80 1606 80 1658
rect 132 1606 170 1658
rect -170 1441 170 1606
rect -170 1389 -132 1441
rect -80 1389 80 1441
rect 132 1389 170 1441
rect -170 1223 170 1389
rect -170 1171 -132 1223
rect -80 1171 80 1223
rect 132 1171 170 1223
rect -170 1005 170 1171
rect -170 953 -132 1005
rect -80 953 80 1005
rect 132 953 170 1005
rect -170 788 170 953
rect -170 736 -132 788
rect -80 736 80 788
rect 132 736 170 788
rect -170 570 170 736
rect -170 518 -132 570
rect -80 518 80 570
rect 132 518 170 570
rect -170 353 170 518
rect -170 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -170 135 170 301
rect -170 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -170 -83 170 83
rect -170 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -170 -301 170 -135
rect -170 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -170 -518 170 -353
rect -170 -570 -132 -518
rect -80 -570 80 -518
rect 132 -570 170 -518
rect -170 -736 170 -570
rect -170 -788 -132 -736
rect -80 -788 80 -736
rect 132 -788 170 -736
rect -170 -953 170 -788
rect -170 -1005 -132 -953
rect -80 -1005 80 -953
rect 132 -1005 170 -953
rect -170 -1171 170 -1005
rect -170 -1223 -132 -1171
rect -80 -1223 80 -1171
rect 132 -1223 170 -1171
rect -170 -1389 170 -1223
rect -170 -1441 -132 -1389
rect -80 -1441 80 -1389
rect 132 -1441 170 -1389
rect -170 -1606 170 -1441
rect -170 -1658 -132 -1606
rect -80 -1658 80 -1606
rect 132 -1658 170 -1606
rect -170 -1824 170 -1658
rect -170 -1876 -132 -1824
rect -80 -1876 80 -1824
rect 132 -1876 170 -1824
rect -170 -2042 170 -1876
rect -170 -2094 -132 -2042
rect -80 -2094 80 -2042
rect 132 -2094 170 -2042
rect -170 -2259 170 -2094
rect -170 -2311 -132 -2259
rect -80 -2311 80 -2259
rect 132 -2311 170 -2259
rect -170 -2477 170 -2311
rect -170 -2529 -132 -2477
rect -80 -2529 80 -2477
rect 132 -2529 170 -2477
rect -170 -2694 170 -2529
rect -170 -2746 -132 -2694
rect -80 -2746 80 -2694
rect 132 -2746 170 -2694
rect -170 -2912 170 -2746
rect -170 -2964 -132 -2912
rect -80 -2964 80 -2912
rect 132 -2964 170 -2912
rect -170 -3130 170 -2964
rect -170 -3182 -132 -3130
rect -80 -3182 80 -3130
rect 132 -3182 170 -3130
rect -170 -3347 170 -3182
rect -170 -3399 -132 -3347
rect -80 -3399 80 -3347
rect 132 -3399 170 -3347
rect -170 -3565 170 -3399
rect -170 -3617 -132 -3565
rect -80 -3617 80 -3565
rect 132 -3617 170 -3565
rect -170 -3783 170 -3617
rect -170 -3835 -132 -3783
rect -80 -3835 80 -3783
rect 132 -3835 170 -3783
rect -170 -4000 170 -3835
rect -170 -4052 -132 -4000
rect -80 -4052 80 -4000
rect 132 -4052 170 -4000
rect -170 -4218 170 -4052
rect -170 -4270 -132 -4218
rect -80 -4270 80 -4218
rect 132 -4270 170 -4218
rect -170 -4436 170 -4270
rect -170 -4488 -132 -4436
rect -80 -4488 80 -4436
rect 132 -4488 170 -4436
rect -170 -4653 170 -4488
rect -170 -4705 -132 -4653
rect -80 -4705 80 -4653
rect 132 -4705 170 -4653
rect -170 -4871 170 -4705
rect -170 -4923 -132 -4871
rect -80 -4923 80 -4871
rect 132 -4923 170 -4871
rect -170 -5088 170 -4923
rect -170 -5140 -132 -5088
rect -80 -5140 80 -5088
rect 132 -5140 170 -5088
rect -170 -5306 170 -5140
rect -170 -5358 -132 -5306
rect -80 -5358 80 -5306
rect 132 -5358 170 -5306
rect -170 -5524 170 -5358
rect -170 -5576 -132 -5524
rect -80 -5576 80 -5524
rect 132 -5576 170 -5524
rect -170 -5741 170 -5576
rect -170 -5793 -132 -5741
rect -80 -5793 80 -5741
rect 132 -5793 170 -5741
rect -170 -5959 170 -5793
rect -170 -6011 -132 -5959
rect -80 -6011 80 -5959
rect 132 -6011 170 -5959
rect -170 -6177 170 -6011
rect -170 -6229 -132 -6177
rect -80 -6229 80 -6177
rect 132 -6229 170 -6177
rect -170 -6394 170 -6229
rect -170 -6446 -132 -6394
rect -80 -6446 80 -6394
rect 132 -6446 170 -6394
rect -170 -6612 170 -6446
rect -170 -6664 -132 -6612
rect -80 -6664 80 -6612
rect 132 -6664 170 -6612
rect -170 -6829 170 -6664
rect -170 -6881 -132 -6829
rect -80 -6881 80 -6829
rect 132 -6881 170 -6829
rect -170 -7047 170 -6881
rect -170 -7099 -132 -7047
rect -80 -7099 80 -7047
rect 132 -7099 170 -7047
rect -170 -7265 170 -7099
rect -170 -7317 -132 -7265
rect -80 -7317 80 -7265
rect 132 -7317 170 -7265
rect -170 -7482 170 -7317
rect -170 -7534 -132 -7482
rect -80 -7534 80 -7482
rect 132 -7534 170 -7482
rect -170 -7700 170 -7534
rect -170 -7752 -132 -7700
rect -80 -7752 80 -7700
rect 132 -7752 170 -7700
rect -170 -7918 170 -7752
rect -170 -7970 -132 -7918
rect -80 -7970 80 -7918
rect 132 -7970 170 -7918
rect -170 -8135 170 -7970
rect -170 -8187 -132 -8135
rect -80 -8187 80 -8135
rect 132 -8187 170 -8135
rect -170 -8353 170 -8187
rect -170 -8405 -132 -8353
rect -80 -8405 80 -8353
rect 132 -8405 170 -8353
rect -170 -8571 170 -8405
rect -170 -8623 -132 -8571
rect -80 -8623 80 -8571
rect 132 -8623 170 -8571
rect -170 -8788 170 -8623
rect -170 -8840 -132 -8788
rect -80 -8840 80 -8788
rect 132 -8840 170 -8788
rect -170 -9006 170 -8840
rect -170 -9058 -132 -9006
rect -80 -9058 80 -9006
rect 132 -9058 170 -9006
rect -170 -9223 170 -9058
rect -170 -9275 -132 -9223
rect -80 -9275 80 -9223
rect 132 -9275 170 -9223
rect -170 -9441 170 -9275
rect -170 -9493 -132 -9441
rect -80 -9493 80 -9441
rect 132 -9493 170 -9441
rect -170 -9659 170 -9493
rect -170 -9711 -132 -9659
rect -80 -9711 80 -9659
rect 132 -9711 170 -9659
rect -170 -9876 170 -9711
rect -170 -9928 -132 -9876
rect -80 -9928 80 -9876
rect 132 -9928 170 -9876
rect -170 -10094 170 -9928
rect -170 -10146 -132 -10094
rect -80 -10146 80 -10094
rect 132 -10146 170 -10094
rect -170 -10312 170 -10146
rect -170 -10364 -132 -10312
rect -80 -10364 80 -10312
rect 132 -10364 170 -10312
rect -170 -10529 170 -10364
rect -170 -10581 -132 -10529
rect -80 -10581 80 -10529
rect 132 -10581 170 -10529
rect -170 -10747 170 -10581
rect -170 -10799 -132 -10747
rect -80 -10799 80 -10747
rect 132 -10799 170 -10747
rect -170 -10965 170 -10799
rect -170 -11017 -132 -10965
rect -80 -11017 80 -10965
rect 132 -11017 170 -10965
rect -170 -11182 170 -11017
rect -170 -11234 -132 -11182
rect -80 -11234 80 -11182
rect 132 -11234 170 -11182
rect -170 -11400 170 -11234
rect -170 -11452 -132 -11400
rect -80 -11452 80 -11400
rect 132 -11452 170 -11400
rect -170 -11617 170 -11452
rect -170 -11669 -132 -11617
rect -80 -11669 80 -11617
rect 132 -11669 170 -11617
rect -170 -11835 170 -11669
rect -170 -11887 -132 -11835
rect -80 -11887 80 -11835
rect 132 -11887 170 -11835
rect -170 -12053 170 -11887
rect -170 -12105 -132 -12053
rect -80 -12105 80 -12053
rect 132 -12105 170 -12053
rect -170 -12270 170 -12105
rect -170 -12322 -132 -12270
rect -80 -12322 80 -12270
rect 132 -12322 170 -12270
rect -170 -12488 170 -12322
rect -170 -12540 -132 -12488
rect -80 -12540 80 -12488
rect 132 -12540 170 -12488
rect -170 -12706 170 -12540
rect -170 -12758 -132 -12706
rect -80 -12758 80 -12706
rect 132 -12758 170 -12706
rect -170 -12923 170 -12758
rect -170 -12975 -132 -12923
rect -80 -12975 80 -12923
rect 132 -12975 170 -12923
rect -170 -13141 170 -12975
rect -170 -13193 -132 -13141
rect -80 -13193 80 -13141
rect 132 -13193 170 -13141
rect -170 -13358 170 -13193
rect -170 -13410 -132 -13358
rect -80 -13410 80 -13358
rect 132 -13410 170 -13358
rect -170 -13576 170 -13410
rect -170 -13628 -132 -13576
rect -80 -13628 80 -13576
rect 132 -13628 170 -13576
rect -170 -13794 170 -13628
rect -170 -13846 -132 -13794
rect -80 -13846 80 -13794
rect 132 -13846 170 -13794
rect -170 -14011 170 -13846
rect -170 -14063 -132 -14011
rect -80 -14063 80 -14011
rect 132 -14063 170 -14011
rect -170 -14104 170 -14063
<< via1 >>
rect -132 14011 -80 14063
rect 80 14011 132 14063
rect -132 13794 -80 13846
rect 80 13794 132 13846
rect -132 13576 -80 13628
rect 80 13576 132 13628
rect -132 13358 -80 13410
rect 80 13358 132 13410
rect -132 13141 -80 13193
rect 80 13141 132 13193
rect -132 12923 -80 12975
rect 80 12923 132 12975
rect -132 12706 -80 12758
rect 80 12706 132 12758
rect -132 12488 -80 12540
rect 80 12488 132 12540
rect -132 12270 -80 12322
rect 80 12270 132 12322
rect -132 12053 -80 12105
rect 80 12053 132 12105
rect -132 11835 -80 11887
rect 80 11835 132 11887
rect -132 11617 -80 11669
rect 80 11617 132 11669
rect -132 11400 -80 11452
rect 80 11400 132 11452
rect -132 11182 -80 11234
rect 80 11182 132 11234
rect -132 10965 -80 11017
rect 80 10965 132 11017
rect -132 10747 -80 10799
rect 80 10747 132 10799
rect -132 10529 -80 10581
rect 80 10529 132 10581
rect -132 10312 -80 10364
rect 80 10312 132 10364
rect -132 10094 -80 10146
rect 80 10094 132 10146
rect -132 9876 -80 9928
rect 80 9876 132 9928
rect -132 9659 -80 9711
rect 80 9659 132 9711
rect -132 9441 -80 9493
rect 80 9441 132 9493
rect -132 9223 -80 9275
rect 80 9223 132 9275
rect -132 9006 -80 9058
rect 80 9006 132 9058
rect -132 8788 -80 8840
rect 80 8788 132 8840
rect -132 8571 -80 8623
rect 80 8571 132 8623
rect -132 8353 -80 8405
rect 80 8353 132 8405
rect -132 8135 -80 8187
rect 80 8135 132 8187
rect -132 7918 -80 7970
rect 80 7918 132 7970
rect -132 7700 -80 7752
rect 80 7700 132 7752
rect -132 7482 -80 7534
rect 80 7482 132 7534
rect -132 7265 -80 7317
rect 80 7265 132 7317
rect -132 7047 -80 7099
rect 80 7047 132 7099
rect -132 6829 -80 6881
rect 80 6829 132 6881
rect -132 6612 -80 6664
rect 80 6612 132 6664
rect -132 6394 -80 6446
rect 80 6394 132 6446
rect -132 6177 -80 6229
rect 80 6177 132 6229
rect -132 5959 -80 6011
rect 80 5959 132 6011
rect -132 5741 -80 5793
rect 80 5741 132 5793
rect -132 5524 -80 5576
rect 80 5524 132 5576
rect -132 5306 -80 5358
rect 80 5306 132 5358
rect -132 5088 -80 5140
rect 80 5088 132 5140
rect -132 4871 -80 4923
rect 80 4871 132 4923
rect -132 4653 -80 4705
rect 80 4653 132 4705
rect -132 4436 -80 4488
rect 80 4436 132 4488
rect -132 4218 -80 4270
rect 80 4218 132 4270
rect -132 4000 -80 4052
rect 80 4000 132 4052
rect -132 3783 -80 3835
rect 80 3783 132 3835
rect -132 3565 -80 3617
rect 80 3565 132 3617
rect -132 3347 -80 3399
rect 80 3347 132 3399
rect -132 3130 -80 3182
rect 80 3130 132 3182
rect -132 2912 -80 2964
rect 80 2912 132 2964
rect -132 2694 -80 2746
rect 80 2694 132 2746
rect -132 2477 -80 2529
rect 80 2477 132 2529
rect -132 2259 -80 2311
rect 80 2259 132 2311
rect -132 2042 -80 2094
rect 80 2042 132 2094
rect -132 1824 -80 1876
rect 80 1824 132 1876
rect -132 1606 -80 1658
rect 80 1606 132 1658
rect -132 1389 -80 1441
rect 80 1389 132 1441
rect -132 1171 -80 1223
rect 80 1171 132 1223
rect -132 953 -80 1005
rect 80 953 132 1005
rect -132 736 -80 788
rect 80 736 132 788
rect -132 518 -80 570
rect 80 518 132 570
rect -132 301 -80 353
rect 80 301 132 353
rect -132 83 -80 135
rect 80 83 132 135
rect -132 -135 -80 -83
rect 80 -135 132 -83
rect -132 -353 -80 -301
rect 80 -353 132 -301
rect -132 -570 -80 -518
rect 80 -570 132 -518
rect -132 -788 -80 -736
rect 80 -788 132 -736
rect -132 -1005 -80 -953
rect 80 -1005 132 -953
rect -132 -1223 -80 -1171
rect 80 -1223 132 -1171
rect -132 -1441 -80 -1389
rect 80 -1441 132 -1389
rect -132 -1658 -80 -1606
rect 80 -1658 132 -1606
rect -132 -1876 -80 -1824
rect 80 -1876 132 -1824
rect -132 -2094 -80 -2042
rect 80 -2094 132 -2042
rect -132 -2311 -80 -2259
rect 80 -2311 132 -2259
rect -132 -2529 -80 -2477
rect 80 -2529 132 -2477
rect -132 -2746 -80 -2694
rect 80 -2746 132 -2694
rect -132 -2964 -80 -2912
rect 80 -2964 132 -2912
rect -132 -3182 -80 -3130
rect 80 -3182 132 -3130
rect -132 -3399 -80 -3347
rect 80 -3399 132 -3347
rect -132 -3617 -80 -3565
rect 80 -3617 132 -3565
rect -132 -3835 -80 -3783
rect 80 -3835 132 -3783
rect -132 -4052 -80 -4000
rect 80 -4052 132 -4000
rect -132 -4270 -80 -4218
rect 80 -4270 132 -4218
rect -132 -4488 -80 -4436
rect 80 -4488 132 -4436
rect -132 -4705 -80 -4653
rect 80 -4705 132 -4653
rect -132 -4923 -80 -4871
rect 80 -4923 132 -4871
rect -132 -5140 -80 -5088
rect 80 -5140 132 -5088
rect -132 -5358 -80 -5306
rect 80 -5358 132 -5306
rect -132 -5576 -80 -5524
rect 80 -5576 132 -5524
rect -132 -5793 -80 -5741
rect 80 -5793 132 -5741
rect -132 -6011 -80 -5959
rect 80 -6011 132 -5959
rect -132 -6229 -80 -6177
rect 80 -6229 132 -6177
rect -132 -6446 -80 -6394
rect 80 -6446 132 -6394
rect -132 -6664 -80 -6612
rect 80 -6664 132 -6612
rect -132 -6881 -80 -6829
rect 80 -6881 132 -6829
rect -132 -7099 -80 -7047
rect 80 -7099 132 -7047
rect -132 -7317 -80 -7265
rect 80 -7317 132 -7265
rect -132 -7534 -80 -7482
rect 80 -7534 132 -7482
rect -132 -7752 -80 -7700
rect 80 -7752 132 -7700
rect -132 -7970 -80 -7918
rect 80 -7970 132 -7918
rect -132 -8187 -80 -8135
rect 80 -8187 132 -8135
rect -132 -8405 -80 -8353
rect 80 -8405 132 -8353
rect -132 -8623 -80 -8571
rect 80 -8623 132 -8571
rect -132 -8840 -80 -8788
rect 80 -8840 132 -8788
rect -132 -9058 -80 -9006
rect 80 -9058 132 -9006
rect -132 -9275 -80 -9223
rect 80 -9275 132 -9223
rect -132 -9493 -80 -9441
rect 80 -9493 132 -9441
rect -132 -9711 -80 -9659
rect 80 -9711 132 -9659
rect -132 -9928 -80 -9876
rect 80 -9928 132 -9876
rect -132 -10146 -80 -10094
rect 80 -10146 132 -10094
rect -132 -10364 -80 -10312
rect 80 -10364 132 -10312
rect -132 -10581 -80 -10529
rect 80 -10581 132 -10529
rect -132 -10799 -80 -10747
rect 80 -10799 132 -10747
rect -132 -11017 -80 -10965
rect 80 -11017 132 -10965
rect -132 -11234 -80 -11182
rect 80 -11234 132 -11182
rect -132 -11452 -80 -11400
rect 80 -11452 132 -11400
rect -132 -11669 -80 -11617
rect 80 -11669 132 -11617
rect -132 -11887 -80 -11835
rect 80 -11887 132 -11835
rect -132 -12105 -80 -12053
rect 80 -12105 132 -12053
rect -132 -12322 -80 -12270
rect 80 -12322 132 -12270
rect -132 -12540 -80 -12488
rect 80 -12540 132 -12488
rect -132 -12758 -80 -12706
rect 80 -12758 132 -12706
rect -132 -12975 -80 -12923
rect 80 -12975 132 -12923
rect -132 -13193 -80 -13141
rect 80 -13193 132 -13141
rect -132 -13410 -80 -13358
rect 80 -13410 132 -13358
rect -132 -13628 -80 -13576
rect 80 -13628 132 -13576
rect -132 -13846 -80 -13794
rect 80 -13846 132 -13794
rect -132 -14063 -80 -14011
rect 80 -14063 132 -14011
<< metal2 >>
rect -170 14063 170 14104
rect -170 14011 -132 14063
rect -80 14011 80 14063
rect 132 14011 170 14063
rect -170 13846 170 14011
rect -170 13794 -132 13846
rect -80 13794 80 13846
rect 132 13794 170 13846
rect -170 13628 170 13794
rect -170 13576 -132 13628
rect -80 13576 80 13628
rect 132 13576 170 13628
rect -170 13410 170 13576
rect -170 13358 -132 13410
rect -80 13358 80 13410
rect 132 13358 170 13410
rect -170 13193 170 13358
rect -170 13141 -132 13193
rect -80 13141 80 13193
rect 132 13141 170 13193
rect -170 12975 170 13141
rect -170 12923 -132 12975
rect -80 12923 80 12975
rect 132 12923 170 12975
rect -170 12758 170 12923
rect -170 12706 -132 12758
rect -80 12706 80 12758
rect 132 12706 170 12758
rect -170 12540 170 12706
rect -170 12488 -132 12540
rect -80 12488 80 12540
rect 132 12488 170 12540
rect -170 12322 170 12488
rect -170 12270 -132 12322
rect -80 12270 80 12322
rect 132 12270 170 12322
rect -170 12105 170 12270
rect -170 12053 -132 12105
rect -80 12053 80 12105
rect 132 12053 170 12105
rect -170 11887 170 12053
rect -170 11835 -132 11887
rect -80 11835 80 11887
rect 132 11835 170 11887
rect -170 11669 170 11835
rect -170 11617 -132 11669
rect -80 11617 80 11669
rect 132 11617 170 11669
rect -170 11452 170 11617
rect -170 11400 -132 11452
rect -80 11400 80 11452
rect 132 11400 170 11452
rect -170 11234 170 11400
rect -170 11182 -132 11234
rect -80 11182 80 11234
rect 132 11182 170 11234
rect -170 11017 170 11182
rect -170 10965 -132 11017
rect -80 10965 80 11017
rect 132 10965 170 11017
rect -170 10799 170 10965
rect -170 10747 -132 10799
rect -80 10747 80 10799
rect 132 10747 170 10799
rect -170 10581 170 10747
rect -170 10529 -132 10581
rect -80 10529 80 10581
rect 132 10529 170 10581
rect -170 10364 170 10529
rect -170 10312 -132 10364
rect -80 10312 80 10364
rect 132 10312 170 10364
rect -170 10146 170 10312
rect -170 10094 -132 10146
rect -80 10094 80 10146
rect 132 10094 170 10146
rect -170 9928 170 10094
rect -170 9876 -132 9928
rect -80 9876 80 9928
rect 132 9876 170 9928
rect -170 9711 170 9876
rect -170 9659 -132 9711
rect -80 9659 80 9711
rect 132 9659 170 9711
rect -170 9493 170 9659
rect -170 9441 -132 9493
rect -80 9441 80 9493
rect 132 9441 170 9493
rect -170 9275 170 9441
rect -170 9223 -132 9275
rect -80 9223 80 9275
rect 132 9223 170 9275
rect -170 9058 170 9223
rect -170 9006 -132 9058
rect -80 9006 80 9058
rect 132 9006 170 9058
rect -170 8840 170 9006
rect -170 8788 -132 8840
rect -80 8788 80 8840
rect 132 8788 170 8840
rect -170 8623 170 8788
rect -170 8571 -132 8623
rect -80 8571 80 8623
rect 132 8571 170 8623
rect -170 8405 170 8571
rect -170 8353 -132 8405
rect -80 8353 80 8405
rect 132 8353 170 8405
rect -170 8187 170 8353
rect -170 8135 -132 8187
rect -80 8135 80 8187
rect 132 8135 170 8187
rect -170 7970 170 8135
rect -170 7918 -132 7970
rect -80 7918 80 7970
rect 132 7918 170 7970
rect -170 7752 170 7918
rect -170 7700 -132 7752
rect -80 7700 80 7752
rect 132 7700 170 7752
rect -170 7534 170 7700
rect -170 7482 -132 7534
rect -80 7482 80 7534
rect 132 7482 170 7534
rect -170 7317 170 7482
rect -170 7265 -132 7317
rect -80 7265 80 7317
rect 132 7265 170 7317
rect -170 7099 170 7265
rect -170 7047 -132 7099
rect -80 7047 80 7099
rect 132 7047 170 7099
rect -170 6881 170 7047
rect -170 6829 -132 6881
rect -80 6829 80 6881
rect 132 6829 170 6881
rect -170 6664 170 6829
rect -170 6612 -132 6664
rect -80 6612 80 6664
rect 132 6612 170 6664
rect -170 6446 170 6612
rect -170 6394 -132 6446
rect -80 6394 80 6446
rect 132 6394 170 6446
rect -170 6229 170 6394
rect -170 6177 -132 6229
rect -80 6177 80 6229
rect 132 6177 170 6229
rect -170 6011 170 6177
rect -170 5959 -132 6011
rect -80 5959 80 6011
rect 132 5959 170 6011
rect -170 5793 170 5959
rect -170 5741 -132 5793
rect -80 5741 80 5793
rect 132 5741 170 5793
rect -170 5576 170 5741
rect -170 5524 -132 5576
rect -80 5524 80 5576
rect 132 5524 170 5576
rect -170 5358 170 5524
rect -170 5306 -132 5358
rect -80 5306 80 5358
rect 132 5306 170 5358
rect -170 5140 170 5306
rect -170 5088 -132 5140
rect -80 5088 80 5140
rect 132 5088 170 5140
rect -170 4923 170 5088
rect -170 4871 -132 4923
rect -80 4871 80 4923
rect 132 4871 170 4923
rect -170 4705 170 4871
rect -170 4653 -132 4705
rect -80 4653 80 4705
rect 132 4653 170 4705
rect -170 4488 170 4653
rect -170 4436 -132 4488
rect -80 4436 80 4488
rect 132 4436 170 4488
rect -170 4270 170 4436
rect -170 4218 -132 4270
rect -80 4218 80 4270
rect 132 4218 170 4270
rect -170 4052 170 4218
rect -170 4000 -132 4052
rect -80 4000 80 4052
rect 132 4000 170 4052
rect -170 3835 170 4000
rect -170 3783 -132 3835
rect -80 3783 80 3835
rect 132 3783 170 3835
rect -170 3617 170 3783
rect -170 3565 -132 3617
rect -80 3565 80 3617
rect 132 3565 170 3617
rect -170 3399 170 3565
rect -170 3347 -132 3399
rect -80 3347 80 3399
rect 132 3347 170 3399
rect -170 3182 170 3347
rect -170 3130 -132 3182
rect -80 3130 80 3182
rect 132 3130 170 3182
rect -170 2964 170 3130
rect -170 2912 -132 2964
rect -80 2912 80 2964
rect 132 2912 170 2964
rect -170 2746 170 2912
rect -170 2694 -132 2746
rect -80 2694 80 2746
rect 132 2694 170 2746
rect -170 2529 170 2694
rect -170 2477 -132 2529
rect -80 2477 80 2529
rect 132 2477 170 2529
rect -170 2311 170 2477
rect -170 2259 -132 2311
rect -80 2259 80 2311
rect 132 2259 170 2311
rect -170 2094 170 2259
rect -170 2042 -132 2094
rect -80 2042 80 2094
rect 132 2042 170 2094
rect -170 1876 170 2042
rect -170 1824 -132 1876
rect -80 1824 80 1876
rect 132 1824 170 1876
rect -170 1658 170 1824
rect -170 1606 -132 1658
rect -80 1606 80 1658
rect 132 1606 170 1658
rect -170 1441 170 1606
rect -170 1389 -132 1441
rect -80 1389 80 1441
rect 132 1389 170 1441
rect -170 1223 170 1389
rect -170 1171 -132 1223
rect -80 1171 80 1223
rect 132 1171 170 1223
rect -170 1005 170 1171
rect -170 953 -132 1005
rect -80 953 80 1005
rect 132 953 170 1005
rect -170 788 170 953
rect -170 736 -132 788
rect -80 736 80 788
rect 132 736 170 788
rect -170 570 170 736
rect -170 518 -132 570
rect -80 518 80 570
rect 132 518 170 570
rect -170 353 170 518
rect -170 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -170 135 170 301
rect -170 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -170 -83 170 83
rect -170 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -170 -301 170 -135
rect -170 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -170 -518 170 -353
rect -170 -570 -132 -518
rect -80 -570 80 -518
rect 132 -570 170 -518
rect -170 -736 170 -570
rect -170 -788 -132 -736
rect -80 -788 80 -736
rect 132 -788 170 -736
rect -170 -953 170 -788
rect -170 -1005 -132 -953
rect -80 -1005 80 -953
rect 132 -1005 170 -953
rect -170 -1171 170 -1005
rect -170 -1223 -132 -1171
rect -80 -1223 80 -1171
rect 132 -1223 170 -1171
rect -170 -1389 170 -1223
rect -170 -1441 -132 -1389
rect -80 -1441 80 -1389
rect 132 -1441 170 -1389
rect -170 -1606 170 -1441
rect -170 -1658 -132 -1606
rect -80 -1658 80 -1606
rect 132 -1658 170 -1606
rect -170 -1824 170 -1658
rect -170 -1876 -132 -1824
rect -80 -1876 80 -1824
rect 132 -1876 170 -1824
rect -170 -2042 170 -1876
rect -170 -2094 -132 -2042
rect -80 -2094 80 -2042
rect 132 -2094 170 -2042
rect -170 -2259 170 -2094
rect -170 -2311 -132 -2259
rect -80 -2311 80 -2259
rect 132 -2311 170 -2259
rect -170 -2477 170 -2311
rect -170 -2529 -132 -2477
rect -80 -2529 80 -2477
rect 132 -2529 170 -2477
rect -170 -2694 170 -2529
rect -170 -2746 -132 -2694
rect -80 -2746 80 -2694
rect 132 -2746 170 -2694
rect -170 -2912 170 -2746
rect -170 -2964 -132 -2912
rect -80 -2964 80 -2912
rect 132 -2964 170 -2912
rect -170 -3130 170 -2964
rect -170 -3182 -132 -3130
rect -80 -3182 80 -3130
rect 132 -3182 170 -3130
rect -170 -3347 170 -3182
rect -170 -3399 -132 -3347
rect -80 -3399 80 -3347
rect 132 -3399 170 -3347
rect -170 -3565 170 -3399
rect -170 -3617 -132 -3565
rect -80 -3617 80 -3565
rect 132 -3617 170 -3565
rect -170 -3783 170 -3617
rect -170 -3835 -132 -3783
rect -80 -3835 80 -3783
rect 132 -3835 170 -3783
rect -170 -4000 170 -3835
rect -170 -4052 -132 -4000
rect -80 -4052 80 -4000
rect 132 -4052 170 -4000
rect -170 -4218 170 -4052
rect -170 -4270 -132 -4218
rect -80 -4270 80 -4218
rect 132 -4270 170 -4218
rect -170 -4436 170 -4270
rect -170 -4488 -132 -4436
rect -80 -4488 80 -4436
rect 132 -4488 170 -4436
rect -170 -4653 170 -4488
rect -170 -4705 -132 -4653
rect -80 -4705 80 -4653
rect 132 -4705 170 -4653
rect -170 -4871 170 -4705
rect -170 -4923 -132 -4871
rect -80 -4923 80 -4871
rect 132 -4923 170 -4871
rect -170 -5088 170 -4923
rect -170 -5140 -132 -5088
rect -80 -5140 80 -5088
rect 132 -5140 170 -5088
rect -170 -5306 170 -5140
rect -170 -5358 -132 -5306
rect -80 -5358 80 -5306
rect 132 -5358 170 -5306
rect -170 -5524 170 -5358
rect -170 -5576 -132 -5524
rect -80 -5576 80 -5524
rect 132 -5576 170 -5524
rect -170 -5741 170 -5576
rect -170 -5793 -132 -5741
rect -80 -5793 80 -5741
rect 132 -5793 170 -5741
rect -170 -5959 170 -5793
rect -170 -6011 -132 -5959
rect -80 -6011 80 -5959
rect 132 -6011 170 -5959
rect -170 -6177 170 -6011
rect -170 -6229 -132 -6177
rect -80 -6229 80 -6177
rect 132 -6229 170 -6177
rect -170 -6394 170 -6229
rect -170 -6446 -132 -6394
rect -80 -6446 80 -6394
rect 132 -6446 170 -6394
rect -170 -6612 170 -6446
rect -170 -6664 -132 -6612
rect -80 -6664 80 -6612
rect 132 -6664 170 -6612
rect -170 -6829 170 -6664
rect -170 -6881 -132 -6829
rect -80 -6881 80 -6829
rect 132 -6881 170 -6829
rect -170 -7047 170 -6881
rect -170 -7099 -132 -7047
rect -80 -7099 80 -7047
rect 132 -7099 170 -7047
rect -170 -7265 170 -7099
rect -170 -7317 -132 -7265
rect -80 -7317 80 -7265
rect 132 -7317 170 -7265
rect -170 -7482 170 -7317
rect -170 -7534 -132 -7482
rect -80 -7534 80 -7482
rect 132 -7534 170 -7482
rect -170 -7700 170 -7534
rect -170 -7752 -132 -7700
rect -80 -7752 80 -7700
rect 132 -7752 170 -7700
rect -170 -7918 170 -7752
rect -170 -7970 -132 -7918
rect -80 -7970 80 -7918
rect 132 -7970 170 -7918
rect -170 -8135 170 -7970
rect -170 -8187 -132 -8135
rect -80 -8187 80 -8135
rect 132 -8187 170 -8135
rect -170 -8353 170 -8187
rect -170 -8405 -132 -8353
rect -80 -8405 80 -8353
rect 132 -8405 170 -8353
rect -170 -8571 170 -8405
rect -170 -8623 -132 -8571
rect -80 -8623 80 -8571
rect 132 -8623 170 -8571
rect -170 -8788 170 -8623
rect -170 -8840 -132 -8788
rect -80 -8840 80 -8788
rect 132 -8840 170 -8788
rect -170 -9006 170 -8840
rect -170 -9058 -132 -9006
rect -80 -9058 80 -9006
rect 132 -9058 170 -9006
rect -170 -9223 170 -9058
rect -170 -9275 -132 -9223
rect -80 -9275 80 -9223
rect 132 -9275 170 -9223
rect -170 -9441 170 -9275
rect -170 -9493 -132 -9441
rect -80 -9493 80 -9441
rect 132 -9493 170 -9441
rect -170 -9659 170 -9493
rect -170 -9711 -132 -9659
rect -80 -9711 80 -9659
rect 132 -9711 170 -9659
rect -170 -9876 170 -9711
rect -170 -9928 -132 -9876
rect -80 -9928 80 -9876
rect 132 -9928 170 -9876
rect -170 -10094 170 -9928
rect -170 -10146 -132 -10094
rect -80 -10146 80 -10094
rect 132 -10146 170 -10094
rect -170 -10312 170 -10146
rect -170 -10364 -132 -10312
rect -80 -10364 80 -10312
rect 132 -10364 170 -10312
rect -170 -10529 170 -10364
rect -170 -10581 -132 -10529
rect -80 -10581 80 -10529
rect 132 -10581 170 -10529
rect -170 -10747 170 -10581
rect -170 -10799 -132 -10747
rect -80 -10799 80 -10747
rect 132 -10799 170 -10747
rect -170 -10965 170 -10799
rect -170 -11017 -132 -10965
rect -80 -11017 80 -10965
rect 132 -11017 170 -10965
rect -170 -11182 170 -11017
rect -170 -11234 -132 -11182
rect -80 -11234 80 -11182
rect 132 -11234 170 -11182
rect -170 -11400 170 -11234
rect -170 -11452 -132 -11400
rect -80 -11452 80 -11400
rect 132 -11452 170 -11400
rect -170 -11617 170 -11452
rect -170 -11669 -132 -11617
rect -80 -11669 80 -11617
rect 132 -11669 170 -11617
rect -170 -11835 170 -11669
rect -170 -11887 -132 -11835
rect -80 -11887 80 -11835
rect 132 -11887 170 -11835
rect -170 -12053 170 -11887
rect -170 -12105 -132 -12053
rect -80 -12105 80 -12053
rect 132 -12105 170 -12053
rect -170 -12270 170 -12105
rect -170 -12322 -132 -12270
rect -80 -12322 80 -12270
rect 132 -12322 170 -12270
rect -170 -12488 170 -12322
rect -170 -12540 -132 -12488
rect -80 -12540 80 -12488
rect 132 -12540 170 -12488
rect -170 -12706 170 -12540
rect -170 -12758 -132 -12706
rect -80 -12758 80 -12706
rect 132 -12758 170 -12706
rect -170 -12923 170 -12758
rect -170 -12975 -132 -12923
rect -80 -12975 80 -12923
rect 132 -12975 170 -12923
rect -170 -13141 170 -12975
rect -170 -13193 -132 -13141
rect -80 -13193 80 -13141
rect 132 -13193 170 -13141
rect -170 -13358 170 -13193
rect -170 -13410 -132 -13358
rect -80 -13410 80 -13358
rect 132 -13410 170 -13358
rect -170 -13576 170 -13410
rect -170 -13628 -132 -13576
rect -80 -13628 80 -13576
rect 132 -13628 170 -13576
rect -170 -13794 170 -13628
rect -170 -13846 -132 -13794
rect -80 -13846 80 -13794
rect 132 -13846 170 -13794
rect -170 -14011 170 -13846
rect -170 -14063 -132 -14011
rect -80 -14063 80 -14011
rect 132 -14063 170 -14011
rect -170 -14104 170 -14063
<< properties >>
string GDS_END 2247866
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2231094
<< end >>
