magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 2203 54557 88011 55557
rect 35945 53519 36945 54557
rect 42135 53477 42444 54557
rect 45745 53475 46606 54557
rect 87011 3345 88011 54557
rect 2203 2345 88011 3345
<< metal2 >>
rect 31407 53974 34809 55039
rect 37049 53974 38336 55039
rect 40506 54039 41539 55039
rect 50710 53974 51911 55039
rect 54147 53974 57559 55039
rect 59830 53974 60272 54994
rect 28693 2345 29135 4295
rect 29308 2345 29750 4295
rect 59216 2345 59658 4835
rect 59830 3295 60272 4295
rect 86587 2345 87587 55029
<< metal3 >>
rect 27079 55231 28079 55839
rect 28493 55039 29493 55839
rect 32631 55039 33631 55839
rect 35945 55231 36945 55839
rect 37336 55039 38336 55839
rect 40506 55039 41506 55839
rect 41803 55231 42803 55839
rect 45634 55231 46634 55839
rect 50822 55039 51822 55839
rect 52386 55231 53386 55839
rect 54490 55039 55490 55839
rect 56183 55039 57183 55839
rect 57911 55231 58911 55839
rect 59468 55039 60468 55839
rect 60712 55231 61712 55839
rect 2203 54039 88293 55039
use M2_M14310590548777_128x8m81  M2_M14310590548777_128x8m81_0
timestamp 1666464484
transform 1 0 59432 0 1 3583
box -162 -1216 162 1216
use M2_M14310590548778_128x8m81  M2_M14310590548778_128x8m81_0
timestamp 1666464484
transform 1 0 60052 0 1 4068
box -162 -224 162 224
use M2_M14310590548778_128x8m81  M2_M14310590548778_128x8m81_1
timestamp 1666464484
transform 1 0 28915 0 1 4068
box -162 -224 162 224
use M2_M14310590548782_128x8m81  M2_M14310590548782_128x8m81_0
timestamp 1666464484
transform 1 0 29524 0 1 3317
box -162 -968 162 968
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_0
timestamp 1666464484
transform 1 0 27590 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_1
timestamp 1666464484
transform 1 0 46119 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_2
timestamp 1666464484
transform 1 0 36446 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_3
timestamp 1666464484
transform 1 0 42288 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_4
timestamp 1666464484
transform 1 0 61197 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_5
timestamp 1666464484
transform 1 0 52871 0 1 55395
box -472 -162 472 162
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_6
timestamp 1666464484
transform 1 0 58396 0 1 55395
box -472 -162 472 162
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_0
timestamp 1666464484
transform 1 0 60052 0 1 3820
box -162 -472 162 472
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_1
timestamp 1666464484
transform 1 0 28915 0 1 3820
box -162 -472 162 472
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_0
timestamp 1666464484
transform 1 0 46119 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_1
timestamp 1666464484
transform 1 0 61197 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_2
timestamp 1666464484
transform 1 0 36446 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_3
timestamp 1666464484
transform 1 0 42288 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_4
timestamp 1666464484
transform 1 0 52871 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_5
timestamp 1666464484
transform 1 0 58396 0 1 55395
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_6
timestamp 1666464484
transform 1 0 27590 0 1 55395
box -472 -162 472 162
use M3_M24310590548779_128x8m81  M3_M24310590548779_128x8m81_0
timestamp 1666464484
transform 1 0 37673 0 1 54522
box -596 -472 596 472
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_0
timestamp 1666464484
transform 1 0 34250 0 1 54541
box -410 -472 410 472
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_1
timestamp 1666464484
transform 1 0 31966 0 1 54541
box -410 -472 410 472
use M3_M24310590548780_128x8m81  M3_M24310590548780_128x8m81_2
timestamp 1666464484
transform 1 0 33115 0 1 54541
box -410 -472 410 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_0
timestamp 1666464484
transform 1 0 56683 0 1 54522
box -472 -472 472 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_1
timestamp 1666464484
transform 1 0 28995 0 1 54536
box -472 -472 472 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_2
timestamp 1666464484
transform 1 0 59968 0 1 54522
box -472 -472 472 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_3
timestamp 1666464484
transform 1 0 51322 0 1 54522
box -472 -472 472 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_4
timestamp 1666464484
transform 1 0 54990 0 1 54522
box -472 -472 472 472
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_5
timestamp 1666464484
transform 1 0 41006 0 1 54522
box -472 -472 472 472
use M3_M24310590548784_128x8m81  M3_M24310590548784_128x8m81_0
timestamp 1666464484
transform 1 0 60052 0 1 4068
box -162 -224 162 224
use M3_M24310590548784_128x8m81  M3_M24310590548784_128x8m81_1
timestamp 1666464484
transform 1 0 28915 0 1 4068
box -162 -224 162 224
use power_route_01_128x8m81  power_route_01_128x8m81_0
timestamp 1666464484
transform -1 0 85469 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_1
timestamp 1666464484
transform -1 0 25893 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_2
timestamp 1666464484
transform 1 0 9233 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_3
timestamp 1666464484
transform 1 0 20033 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_4
timestamp 1666464484
transform 1 0 14633 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_5
timestamp 1666464484
transform 1 0 63409 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_6
timestamp 1666464484
transform 1 0 79609 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_7
timestamp 1666464484
transform 1 0 74209 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_8
timestamp 1666464484
transform 1 0 68809 0 1 53414
box -511 0 1714 2425
use power_route_01_128x8m81  power_route_01_128x8m81_9
timestamp 1666464484
transform 1 0 3833 0 1 53414
box -511 0 1714 2425
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_0
timestamp 1666464484
transform 1 0 -1418 0 1 50689
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_1
timestamp 1666464484
transform 1 0 -1418 0 1 47089
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_2
timestamp 1666464484
transform 1 0 -1418 0 1 48889
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_3
timestamp 1666464484
transform 1 0 -1418 0 1 39889
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_4
timestamp 1666464484
transform 1 0 -1418 0 1 41689
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_5
timestamp 1666464484
transform 1 0 -1418 0 1 45289
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_6
timestamp 1666464484
transform 1 0 -1418 0 1 43489
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_7
timestamp 1666464484
transform 1 0 -1418 0 1 38089
box 3339 -250 30611 1350
use power_route_02_a_128x8m81  power_route_02_a_128x8m81_8
timestamp 1666464484
transform 1 0 -1418 0 1 52489
box 3339 -250 30611 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_0
timestamp 1666464484
transform -1 0 91632 0 1 39889
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_1
timestamp 1666464484
transform -1 0 91632 0 1 41689
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_2
timestamp 1666464484
transform -1 0 91632 0 1 43489
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_3
timestamp 1666464484
transform -1 0 91632 0 1 45289
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_4
timestamp 1666464484
transform -1 0 91632 0 1 47089
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_5
timestamp 1666464484
transform -1 0 91632 0 1 48889
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_6
timestamp 1666464484
transform -1 0 91632 0 1 50689
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_7
timestamp 1666464484
transform -1 0 91632 0 1 52489
box 3339 -250 30290 1350
use power_route_02_b_128x8m81  power_route_02_b_128x8m81_8
timestamp 1666464484
transform -1 0 91632 0 1 38089
box 3339 -250 30290 1350
use power_route_04_128x8m81  power_route_04_128x8m81_0
timestamp 1666464484
transform -1 0 91632 0 1 244
box 3339 2101 6632 52645
use power_route_04_128x8m81  power_route_04_128x8m81_1
timestamp 1666464484
transform 1 0 -1418 0 1 244
box 3339 2101 6632 52645
use power_route_05_128x8m81  power_route_05_128x8m81_0
timestamp 1666464484
transform 1 0 19656 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_1
timestamp 1666464484
transform 1 0 68432 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_2
timestamp 1666464484
transform 1 0 79232 0 1 230
box -8 2115 1235 7462
use power_route_05_128x8m81  power_route_05_128x8m81_3
timestamp 1666464484
transform 1 0 8856 0 1 230
box -8 2115 1235 7462
use power_route_06_128x8m81  power_route_06_128x8m81_0
timestamp 1666464484
transform 1 0 61241 0 1 230
box -7 2115 1234 18431
use power_route_06_128x8m81  power_route_06_128x8m81_1
timestamp 1666464484
transform 1 0 26784 0 1 230
box -7 2115 1234 18431
use power_route_07_128x8m81  power_route_07_128x8m81_0
timestamp 1666464484
transform 1 0 40746 0 1 230
box -8 3065 1235 7462
use power_route_07_128x8m81  power_route_07_128x8m81_1
timestamp 1666464484
transform 1 0 38926 0 1 230
box -8 3065 1235 7462
<< properties >>
string GDS_END 2287216
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2281500
string path 274.950 279.195 274.950 270.195 
<< end >>
