magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 310 1094
<< pwell >>
rect -86 -86 310 453
<< mvpdiode >>
rect 36 632 108 686
rect 36 586 49 632
rect 95 586 108 632
rect 36 573 108 586
<< mvndiode >>
rect 36 320 108 333
rect 36 274 49 320
rect 95 274 108 320
rect 36 220 108 274
<< mvpdiodec >>
rect 49 586 95 632
<< mvndiodec >>
rect 49 274 95 320
<< metal1 >>
rect 0 918 224 1098
rect 30 632 95 643
rect 30 586 49 632
rect 30 320 95 586
rect 30 274 49 320
rect 30 263 95 274
rect 0 -90 224 90
<< labels >>
flabel metal1 s 30 263 95 643 0 FreeSans 200 0 0 0 I
port 1 nsew default input
flabel metal1 s 0 918 224 1098 0 FreeSans 200 0 0 0 VDD
port 2 nsew power bidirectional abutment
flabel metal1 s 0 -90 224 90 0 FreeSans 200 0 0 0 VSS
port 5 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
<< properties >>
string FIXED_BBOX 0 0 224 1008
string GDS_END 1144494
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1143014
string LEFclass core gf180mcu_fd_sc_mcu9t5v0__antennaCELL
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
