magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -697 380 697 393
rect -696 355 697 380
rect -696 299 -661 355
rect -605 299 -450 355
rect -394 299 -239 355
rect -183 299 -28 355
rect 28 299 183 355
rect 239 299 394 355
rect 450 299 605 355
rect 661 299 697 355
rect -696 137 697 299
rect -696 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 697 137
rect -696 -81 697 81
rect -696 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 697 -81
rect -696 -299 697 -137
rect -696 -355 -661 -299
rect -605 -355 -450 -299
rect -394 -355 -239 -299
rect -183 -355 -28 -299
rect 28 -355 183 -299
rect 239 -355 394 -299
rect 450 -355 605 -299
rect 661 -355 697 -299
rect -696 -393 697 -355
<< via2 >>
rect -661 299 -605 355
rect -450 299 -394 355
rect -239 299 -183 355
rect -28 299 28 355
rect 183 299 239 355
rect 394 299 450 355
rect 605 299 661 355
rect -661 81 -605 137
rect -450 81 -394 137
rect -239 81 -183 137
rect -28 81 28 137
rect 183 81 239 137
rect 394 81 450 137
rect 605 81 661 137
rect -661 -137 -605 -81
rect -450 -137 -394 -81
rect -239 -137 -183 -81
rect -28 -137 28 -81
rect 183 -137 239 -81
rect 394 -137 450 -81
rect 605 -137 661 -81
rect -661 -355 -605 -299
rect -450 -355 -394 -299
rect -239 -355 -183 -299
rect -28 -355 28 -299
rect 183 -355 239 -299
rect 394 -355 450 -299
rect 605 -355 661 -299
<< metal3 >>
rect -696 355 697 393
rect -696 299 -661 355
rect -605 299 -450 355
rect -394 299 -239 355
rect -183 299 -28 355
rect 28 299 183 355
rect 239 299 394 355
rect 450 299 605 355
rect 661 299 697 355
rect -696 137 697 299
rect -696 81 -661 137
rect -605 81 -450 137
rect -394 81 -239 137
rect -183 81 -28 137
rect 28 81 183 137
rect 239 81 394 137
rect 450 81 605 137
rect 661 81 697 137
rect -696 -81 697 81
rect -696 -137 -661 -81
rect -605 -137 -450 -81
rect -394 -137 -239 -81
rect -183 -137 -28 -81
rect 28 -137 183 -81
rect 239 -137 394 -81
rect 450 -137 605 -81
rect 661 -137 697 -81
rect -696 -299 697 -137
rect -696 -355 -661 -299
rect -605 -355 -450 -299
rect -394 -355 -239 -299
rect -183 -355 -28 -299
rect 28 -355 183 -299
rect 239 -355 394 -299
rect 450 -355 605 -299
rect 661 -355 697 -299
rect -696 -393 697 -355
<< properties >>
string GDS_END 775124
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 773184
<< end >>
