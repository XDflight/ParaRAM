magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -42 66223 342 66242
rect -42 -23 -23 66223
rect 323 -23 342 66223
rect -42 -42 342 -23
<< psubdiffcont >>
rect -23 -23 323 66223
<< metal1 >>
rect -34 66223 334 66234
rect -34 -23 -23 66223
rect 323 -23 334 66223
rect -34 -34 334 -23
<< properties >>
string GDS_END 1412530
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1242606
<< end >>
