magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 7926 870
rect -86 352 699 377
rect 2089 352 7926 377
<< pwell >>
rect 699 352 2089 377
rect -86 -86 7926 352
<< mvnmos >>
rect 145 68 265 232
rect 369 68 489 232
rect 593 68 713 232
rect 1139 68 1259 232
rect 1451 68 1571 232
rect 1763 68 1883 232
rect 2075 68 2195 232
rect 2387 68 2507 232
rect 2611 68 2731 232
rect 2835 68 2955 232
rect 3059 68 3179 232
rect 3283 68 3403 232
rect 3507 68 3627 232
rect 3767 68 3887 232
rect 3991 68 4111 232
rect 4215 68 4335 232
rect 4439 68 4559 232
rect 4663 68 4783 232
rect 4887 68 5007 232
rect 5111 68 5231 232
rect 5335 68 5455 232
rect 5559 68 5679 232
rect 5783 68 5903 232
rect 6007 68 6127 232
rect 6231 68 6351 232
rect 6455 68 6575 232
rect 6679 68 6799 232
rect 6903 68 7023 232
rect 7127 68 7247 232
rect 7351 68 7471 232
rect 7575 68 7695 232
<< mvpmos >>
rect 208 497 308 716
rect 412 497 512 716
rect 616 497 716 716
rect 1139 497 1239 716
rect 1451 497 1551 716
rect 1763 497 1863 716
rect 2075 497 2175 716
rect 2387 480 2487 716
rect 2611 480 2711 716
rect 2835 480 2935 716
rect 3059 480 3159 716
rect 3283 480 3383 716
rect 3507 480 3607 716
rect 3767 480 3867 716
rect 3991 480 4091 716
rect 4225 480 4325 716
rect 4439 480 4539 716
rect 4663 480 4763 716
rect 4887 480 4987 716
rect 5111 480 5211 716
rect 5335 480 5435 716
rect 5559 480 5659 716
rect 5783 480 5883 716
rect 6007 480 6107 716
rect 6231 480 6331 716
rect 6455 480 6555 716
rect 6679 480 6779 716
rect 6903 480 7003 716
rect 7127 480 7227 716
rect 7351 480 7451 716
rect 7575 480 7675 716
<< mvndiff >>
rect 773 244 845 257
rect 773 232 786 244
rect 57 192 145 232
rect 57 146 70 192
rect 116 146 145 192
rect 57 68 145 146
rect 265 139 369 232
rect 265 93 294 139
rect 340 93 369 139
rect 265 68 369 93
rect 489 166 593 232
rect 489 120 518 166
rect 564 120 593 166
rect 489 68 593 120
rect 713 198 786 232
rect 832 198 845 244
rect 1319 244 1391 257
rect 1319 232 1332 244
rect 713 68 845 198
rect 1007 95 1139 232
rect 1007 49 1020 95
rect 1066 68 1139 95
rect 1259 198 1332 232
rect 1378 232 1391 244
rect 1943 244 2015 257
rect 1943 232 1956 244
rect 1378 198 1451 232
rect 1259 68 1451 198
rect 1571 95 1763 232
rect 1571 68 1644 95
rect 1066 49 1079 68
rect 1007 36 1079 49
rect 1631 49 1644 68
rect 1690 68 1763 95
rect 1883 198 1956 232
rect 2002 232 2015 244
rect 2002 198 2075 232
rect 1883 68 2075 198
rect 2195 95 2387 232
rect 2195 68 2268 95
rect 1690 49 1703 68
rect 1631 36 1703 49
rect 2255 49 2268 68
rect 2314 68 2387 95
rect 2507 192 2611 232
rect 2507 146 2536 192
rect 2582 146 2611 192
rect 2507 68 2611 146
rect 2731 163 2835 232
rect 2731 117 2760 163
rect 2806 117 2835 163
rect 2731 68 2835 117
rect 2955 163 3059 232
rect 2955 117 2984 163
rect 3030 117 3059 163
rect 2955 68 3059 117
rect 3179 163 3283 232
rect 3179 117 3208 163
rect 3254 117 3283 163
rect 3179 68 3283 117
rect 3403 163 3507 232
rect 3403 117 3432 163
rect 3478 117 3507 163
rect 3403 68 3507 117
rect 3627 163 3767 232
rect 3627 117 3656 163
rect 3702 117 3767 163
rect 3627 68 3767 117
rect 3887 163 3991 232
rect 3887 117 3916 163
rect 3962 117 3991 163
rect 3887 68 3991 117
rect 4111 163 4215 232
rect 4111 117 4140 163
rect 4186 117 4215 163
rect 4111 68 4215 117
rect 4335 219 4439 232
rect 4335 173 4364 219
rect 4410 173 4439 219
rect 4335 68 4439 173
rect 4559 127 4663 232
rect 4559 81 4588 127
rect 4634 81 4663 127
rect 4559 68 4663 81
rect 4783 219 4887 232
rect 4783 173 4812 219
rect 4858 173 4887 219
rect 4783 68 4887 173
rect 5007 127 5111 232
rect 5007 81 5036 127
rect 5082 81 5111 127
rect 5007 68 5111 81
rect 5231 219 5335 232
rect 5231 173 5260 219
rect 5306 173 5335 219
rect 5231 68 5335 173
rect 5455 127 5559 232
rect 5455 81 5484 127
rect 5530 81 5559 127
rect 5455 68 5559 81
rect 5679 219 5783 232
rect 5679 173 5708 219
rect 5754 173 5783 219
rect 5679 68 5783 173
rect 5903 127 6007 232
rect 5903 81 5932 127
rect 5978 81 6007 127
rect 5903 68 6007 81
rect 6127 219 6231 232
rect 6127 173 6156 219
rect 6202 173 6231 219
rect 6127 68 6231 173
rect 6351 127 6455 232
rect 6351 81 6380 127
rect 6426 81 6455 127
rect 6351 68 6455 81
rect 6575 219 6679 232
rect 6575 173 6604 219
rect 6650 173 6679 219
rect 6575 68 6679 173
rect 6799 127 6903 232
rect 6799 81 6828 127
rect 6874 81 6903 127
rect 6799 68 6903 81
rect 7023 219 7127 232
rect 7023 173 7052 219
rect 7098 173 7127 219
rect 7023 68 7127 173
rect 7247 127 7351 232
rect 7247 81 7276 127
rect 7322 81 7351 127
rect 7247 68 7351 81
rect 7471 219 7575 232
rect 7471 173 7500 219
rect 7546 173 7575 219
rect 7471 68 7575 173
rect 7695 192 7783 232
rect 7695 146 7724 192
rect 7770 146 7783 192
rect 7695 68 7783 146
rect 2314 49 2327 68
rect 2255 36 2327 49
<< mvpdiff >>
rect 1007 735 1079 748
rect 120 665 208 716
rect 120 525 133 665
rect 179 525 208 665
rect 120 497 208 525
rect 308 703 412 716
rect 308 657 337 703
rect 383 657 412 703
rect 308 497 412 657
rect 512 670 616 716
rect 512 624 541 670
rect 587 624 616 670
rect 512 497 616 624
rect 716 556 804 716
rect 716 510 745 556
rect 791 510 804 556
rect 716 497 804 510
rect 1007 689 1020 735
rect 1066 716 1079 735
rect 1631 735 1703 748
rect 1631 716 1644 735
rect 1066 689 1139 716
rect 1007 497 1139 689
rect 1239 556 1451 716
rect 1239 510 1332 556
rect 1378 510 1451 556
rect 1239 497 1451 510
rect 1551 689 1644 716
rect 1690 716 1703 735
rect 1690 689 1763 716
rect 1551 497 1763 689
rect 1863 556 2075 716
rect 1863 510 1956 556
rect 2002 510 2075 556
rect 1863 497 2075 510
rect 2175 691 2387 716
rect 2175 551 2270 691
rect 2316 551 2387 691
rect 2175 497 2387 551
rect 2239 480 2387 497
rect 2487 665 2611 716
rect 2487 525 2526 665
rect 2572 525 2611 665
rect 2487 480 2611 525
rect 2711 691 2835 716
rect 2711 551 2752 691
rect 2798 551 2835 691
rect 2711 480 2835 551
rect 2935 665 3059 716
rect 2935 525 2976 665
rect 3022 525 3059 665
rect 2935 480 3059 525
rect 3159 691 3283 716
rect 3159 551 3199 691
rect 3245 551 3283 691
rect 3159 480 3283 551
rect 3383 665 3507 716
rect 3383 525 3425 665
rect 3471 525 3507 665
rect 3383 480 3507 525
rect 3607 691 3767 716
rect 3607 551 3666 691
rect 3712 551 3767 691
rect 3607 480 3767 551
rect 3867 665 3991 716
rect 3867 525 3904 665
rect 3950 525 3991 665
rect 3867 480 3991 525
rect 4091 691 4225 716
rect 4091 551 4136 691
rect 4182 551 4225 691
rect 4091 480 4225 551
rect 4325 665 4439 716
rect 4325 525 4364 665
rect 4410 525 4439 665
rect 4325 480 4439 525
rect 4539 703 4663 716
rect 4539 657 4578 703
rect 4624 657 4663 703
rect 4539 480 4663 657
rect 4763 665 4887 716
rect 4763 525 4805 665
rect 4851 525 4887 665
rect 4763 480 4887 525
rect 4987 703 5111 716
rect 4987 657 5027 703
rect 5073 657 5111 703
rect 4987 480 5111 657
rect 5211 665 5335 716
rect 5211 525 5251 665
rect 5297 525 5335 665
rect 5211 480 5335 525
rect 5435 703 5559 716
rect 5435 657 5477 703
rect 5523 657 5559 703
rect 5435 480 5559 657
rect 5659 665 5783 716
rect 5659 525 5702 665
rect 5748 525 5783 665
rect 5659 480 5783 525
rect 5883 703 6007 716
rect 5883 657 5925 703
rect 5971 657 6007 703
rect 5883 480 6007 657
rect 6107 665 6231 716
rect 6107 525 6151 665
rect 6197 525 6231 665
rect 6107 480 6231 525
rect 6331 703 6455 716
rect 6331 657 6373 703
rect 6419 657 6455 703
rect 6331 480 6455 657
rect 6555 665 6679 716
rect 6555 525 6595 665
rect 6641 525 6679 665
rect 6555 480 6679 525
rect 6779 703 6903 716
rect 6779 657 6821 703
rect 6867 657 6903 703
rect 6779 480 6903 657
rect 7003 665 7127 716
rect 7003 525 7045 665
rect 7091 525 7127 665
rect 7003 480 7127 525
rect 7227 703 7351 716
rect 7227 657 7268 703
rect 7314 657 7351 703
rect 7227 480 7351 657
rect 7451 665 7575 716
rect 7451 525 7500 665
rect 7546 525 7575 665
rect 7451 480 7575 525
rect 7675 665 7763 716
rect 7675 525 7704 665
rect 7750 525 7763 665
rect 7675 480 7763 525
<< mvndiffc >>
rect 70 146 116 192
rect 294 93 340 139
rect 518 120 564 166
rect 786 198 832 244
rect 1020 49 1066 95
rect 1332 198 1378 244
rect 1644 49 1690 95
rect 1956 198 2002 244
rect 2268 49 2314 95
rect 2536 146 2582 192
rect 2760 117 2806 163
rect 2984 117 3030 163
rect 3208 117 3254 163
rect 3432 117 3478 163
rect 3656 117 3702 163
rect 3916 117 3962 163
rect 4140 117 4186 163
rect 4364 173 4410 219
rect 4588 81 4634 127
rect 4812 173 4858 219
rect 5036 81 5082 127
rect 5260 173 5306 219
rect 5484 81 5530 127
rect 5708 173 5754 219
rect 5932 81 5978 127
rect 6156 173 6202 219
rect 6380 81 6426 127
rect 6604 173 6650 219
rect 6828 81 6874 127
rect 7052 173 7098 219
rect 7276 81 7322 127
rect 7500 173 7546 219
rect 7724 146 7770 192
<< mvpdiffc >>
rect 133 525 179 665
rect 337 657 383 703
rect 541 624 587 670
rect 745 510 791 556
rect 1020 689 1066 735
rect 1332 510 1378 556
rect 1644 689 1690 735
rect 1956 510 2002 556
rect 2270 551 2316 691
rect 2526 525 2572 665
rect 2752 551 2798 691
rect 2976 525 3022 665
rect 3199 551 3245 691
rect 3425 525 3471 665
rect 3666 551 3712 691
rect 3904 525 3950 665
rect 4136 551 4182 691
rect 4364 525 4410 665
rect 4578 657 4624 703
rect 4805 525 4851 665
rect 5027 657 5073 703
rect 5251 525 5297 665
rect 5477 657 5523 703
rect 5702 525 5748 665
rect 5925 657 5971 703
rect 6151 525 6197 665
rect 6373 657 6419 703
rect 6595 525 6641 665
rect 6821 657 6867 703
rect 7045 525 7091 665
rect 7268 657 7314 703
rect 7500 525 7546 665
rect 7704 525 7750 665
<< polysilicon >>
rect 208 716 308 760
rect 412 716 512 760
rect 616 716 716 760
rect 1139 716 1239 760
rect 1451 716 1551 760
rect 1763 716 1863 760
rect 2075 716 2175 760
rect 2387 716 2487 760
rect 2611 716 2711 760
rect 2835 716 2935 760
rect 3059 716 3159 760
rect 3283 716 3383 760
rect 3507 716 3607 760
rect 3767 716 3867 760
rect 3991 716 4091 760
rect 4225 716 4325 760
rect 4439 716 4539 760
rect 4663 716 4763 760
rect 4887 716 4987 760
rect 5111 716 5211 760
rect 5335 716 5435 760
rect 5559 716 5659 760
rect 5783 716 5883 760
rect 6007 716 6107 760
rect 6231 716 6331 760
rect 6455 716 6555 760
rect 6679 716 6779 760
rect 6903 716 7003 760
rect 7127 716 7227 760
rect 7351 716 7451 760
rect 7575 716 7675 760
rect 208 437 308 497
rect 145 424 308 437
rect 145 378 193 424
rect 239 412 308 424
rect 412 412 512 497
rect 616 464 716 497
rect 616 418 629 464
rect 675 418 716 464
rect 239 378 568 412
rect 616 405 716 418
rect 1139 437 1239 497
rect 1451 437 1551 497
rect 1763 437 1863 497
rect 2075 437 2175 497
rect 1139 424 2175 437
rect 145 372 568 378
rect 145 232 265 372
rect 528 345 568 372
rect 1139 378 1157 424
rect 1959 378 2175 424
rect 1139 365 2175 378
rect 369 311 468 324
rect 369 265 409 311
rect 455 276 468 311
rect 528 305 633 345
rect 593 288 633 305
rect 455 265 489 276
rect 369 232 489 265
rect 593 232 713 288
rect 1139 232 1259 365
rect 145 24 265 68
rect 369 24 489 68
rect 593 24 713 68
rect 1451 232 1571 365
rect 1763 232 1883 365
rect 2075 288 2175 365
rect 2387 399 2487 480
rect 2611 399 2711 480
rect 2835 399 2935 480
rect 3059 399 3159 480
rect 3283 399 3383 480
rect 3507 399 3607 480
rect 3767 399 3867 480
rect 3991 399 4091 480
rect 2387 386 4091 399
rect 2387 340 2406 386
rect 4050 340 4091 386
rect 4225 439 4325 480
rect 4225 393 4249 439
rect 4295 420 4325 439
rect 4439 439 4539 480
rect 4439 420 4467 439
rect 4295 393 4467 420
rect 4513 420 4539 439
rect 4663 439 4763 480
rect 4663 420 4692 439
rect 4513 393 4692 420
rect 4738 420 4763 439
rect 4887 439 4987 480
rect 4887 420 4914 439
rect 4738 393 4914 420
rect 4960 420 4987 439
rect 5111 439 5211 480
rect 5111 420 5139 439
rect 4960 393 5139 420
rect 5185 420 5211 439
rect 5335 439 5435 480
rect 5335 420 5364 439
rect 5185 393 5364 420
rect 5410 420 5435 439
rect 5559 439 5659 480
rect 5559 420 5572 439
rect 5410 393 5572 420
rect 5618 420 5659 439
rect 5783 420 5883 480
rect 6007 420 6107 480
rect 6231 420 6331 480
rect 6455 439 6555 480
rect 6455 420 6482 439
rect 5618 393 6482 420
rect 6528 420 6555 439
rect 6679 439 6779 480
rect 6679 420 6706 439
rect 6528 393 6706 420
rect 6752 420 6779 439
rect 6903 439 7003 480
rect 6903 420 6930 439
rect 6752 393 6930 420
rect 6976 420 7003 439
rect 7127 439 7227 480
rect 7127 420 7153 439
rect 6976 393 7153 420
rect 7199 420 7227 439
rect 7351 439 7451 480
rect 7351 420 7364 439
rect 7199 393 7364 420
rect 7410 420 7451 439
rect 7575 439 7675 480
rect 7575 420 7603 439
rect 7410 393 7603 420
rect 7649 393 7675 439
rect 4225 380 7675 393
rect 2387 327 4091 340
rect 1139 24 1259 68
rect 1451 24 1571 68
rect 2075 232 2195 288
rect 2387 232 2507 327
rect 2611 232 2731 327
rect 2835 232 2955 327
rect 3059 232 3179 327
rect 3283 232 3403 327
rect 3507 232 3627 327
rect 3767 232 3887 327
rect 3991 287 4091 327
rect 4215 319 7695 332
rect 3991 232 4111 287
rect 4215 273 4251 319
rect 4297 292 4479 319
rect 4297 273 4335 292
rect 4215 232 4335 273
rect 4439 273 4479 292
rect 4525 292 4702 319
rect 4525 273 4559 292
rect 4439 232 4559 273
rect 4663 273 4702 292
rect 4748 292 4900 319
rect 4748 273 4783 292
rect 4663 232 4783 273
rect 4887 273 4900 292
rect 4946 292 6964 319
rect 4946 273 5007 292
rect 4887 232 5007 273
rect 5111 232 5231 292
rect 5335 232 5455 292
rect 5559 232 5679 292
rect 5783 232 5903 292
rect 6007 232 6127 292
rect 6231 232 6351 292
rect 6455 232 6575 292
rect 6679 232 6799 292
rect 6903 273 6964 292
rect 7010 292 7163 319
rect 7010 273 7023 292
rect 6903 232 7023 273
rect 7127 273 7163 292
rect 7209 292 7364 319
rect 7209 273 7247 292
rect 7127 232 7247 273
rect 7351 273 7364 292
rect 7410 292 7603 319
rect 7410 273 7471 292
rect 7351 232 7471 273
rect 7575 273 7603 292
rect 7649 273 7695 319
rect 7575 232 7695 273
rect 1763 24 1883 68
rect 2075 24 2195 68
rect 2387 24 2507 68
rect 2611 24 2731 68
rect 2835 24 2955 68
rect 3059 24 3179 68
rect 3283 24 3403 68
rect 3507 24 3627 68
rect 3767 24 3887 68
rect 3991 24 4111 68
rect 4215 24 4335 68
rect 4439 24 4559 68
rect 4663 24 4783 68
rect 4887 24 5007 68
rect 5111 24 5231 68
rect 5335 24 5455 68
rect 5559 24 5679 68
rect 5783 24 5903 68
rect 6007 24 6127 68
rect 6231 24 6351 68
rect 6455 24 6575 68
rect 6679 24 6799 68
rect 6903 24 7023 68
rect 7127 24 7247 68
rect 7351 24 7471 68
rect 7575 24 7695 68
<< polycontact >>
rect 193 378 239 424
rect 629 418 675 464
rect 1157 378 1959 424
rect 409 265 455 311
rect 2406 340 4050 386
rect 4249 393 4295 439
rect 4467 393 4513 439
rect 4692 393 4738 439
rect 4914 393 4960 439
rect 5139 393 5185 439
rect 5364 393 5410 439
rect 5572 393 5618 439
rect 6482 393 6528 439
rect 6706 393 6752 439
rect 6930 393 6976 439
rect 7153 393 7199 439
rect 7364 393 7410 439
rect 7603 393 7649 439
rect 4251 273 4297 319
rect 4479 273 4525 319
rect 4702 273 4748 319
rect 4900 273 4946 319
rect 6964 273 7010 319
rect 7163 273 7209 319
rect 7364 273 7410 319
rect 7603 273 7649 319
<< metal1 >>
rect 0 735 7840 844
rect 0 724 1020 735
rect 326 703 394 724
rect 133 665 179 676
rect 326 657 337 703
rect 383 657 394 703
rect 1009 689 1020 724
rect 1066 724 1644 735
rect 1066 689 1077 724
rect 1631 689 1644 724
rect 1690 724 7840 735
rect 1690 689 1703 724
rect 2270 691 2316 724
rect 518 624 541 670
rect 587 643 963 670
rect 1123 643 1523 671
rect 1771 643 2209 671
rect 587 624 2209 643
rect 837 602 2209 624
rect 837 597 1169 602
rect 1477 597 1817 602
rect 179 525 675 560
rect 133 514 675 525
rect 409 464 675 514
rect 74 424 318 430
rect 74 378 193 424
rect 239 378 318 424
rect 74 354 318 378
rect 409 418 629 464
rect 409 407 675 418
rect 745 556 791 578
rect 409 311 455 407
rect 745 361 791 510
rect 409 245 455 265
rect 70 198 455 245
rect 616 315 791 361
rect 70 192 116 198
rect 616 177 662 315
rect 837 269 883 597
rect 1262 510 1332 556
rect 1378 551 1425 556
rect 1863 551 1956 556
rect 1378 510 1956 551
rect 2002 510 2081 556
rect 1262 505 2081 510
rect 1026 424 1970 430
rect 1026 378 1157 424
rect 1959 378 1970 424
rect 1026 354 1970 378
rect 2035 392 2081 505
rect 2163 485 2209 602
rect 2752 691 2798 724
rect 2270 540 2316 551
rect 2526 665 2572 676
rect 3199 691 3245 724
rect 2752 540 2798 551
rect 2976 665 3022 676
rect 2526 485 2572 525
rect 3666 691 3712 724
rect 3199 540 3245 551
rect 3425 665 3471 676
rect 2976 485 3022 525
rect 4136 691 4182 724
rect 3666 540 3712 551
rect 3904 665 3950 676
rect 3425 485 3471 525
rect 4567 703 4635 724
rect 4136 540 4182 551
rect 4364 665 4410 676
rect 3904 485 3950 525
rect 4567 657 4578 703
rect 4624 657 4635 703
rect 5016 703 5084 724
rect 4805 665 4851 676
rect 4410 525 4805 601
rect 5016 657 5027 703
rect 5073 657 5084 703
rect 5466 703 5534 724
rect 5251 665 5297 676
rect 4851 525 5251 601
rect 5466 657 5477 703
rect 5523 657 5534 703
rect 5914 703 5982 724
rect 5702 665 5748 676
rect 5297 525 5702 601
rect 5914 657 5925 703
rect 5971 657 5982 703
rect 6362 703 6430 724
rect 6151 665 6197 676
rect 5748 525 6151 601
rect 6362 657 6373 703
rect 6419 657 6430 703
rect 6810 703 6878 724
rect 6595 665 6641 676
rect 6197 525 6595 601
rect 6810 657 6821 703
rect 6867 657 6878 703
rect 7257 703 7325 724
rect 7045 665 7091 676
rect 6641 525 7045 601
rect 7257 657 7268 703
rect 7314 657 7325 703
rect 7500 665 7557 676
rect 7091 525 7500 601
rect 7546 525 7557 665
rect 4364 485 7557 525
rect 7704 665 7750 724
rect 7704 506 7750 525
rect 2163 439 4186 485
rect 2163 438 4249 439
rect 4140 393 4249 438
rect 4295 393 4467 439
rect 4513 393 4692 439
rect 4738 393 4914 439
rect 4960 393 5139 439
rect 5185 393 5364 439
rect 5410 393 5572 439
rect 5618 393 5629 439
rect 4140 392 5629 393
rect 2035 386 4065 392
rect 2035 340 2406 386
rect 4050 340 4065 386
rect 2035 326 4065 340
rect 2035 284 2083 326
rect 773 244 883 269
rect 773 198 786 244
rect 832 223 883 244
rect 1319 244 2083 284
rect 4140 273 4251 319
rect 4297 273 4479 319
rect 4525 273 4702 319
rect 4748 273 4900 319
rect 4946 273 4957 319
rect 5790 289 5970 485
rect 6463 393 6482 439
rect 6528 393 6706 439
rect 6752 393 6930 439
rect 6976 393 7153 439
rect 7199 393 7364 439
rect 7410 393 7603 439
rect 7649 393 7660 439
rect 6463 392 7660 393
rect 4140 266 4186 273
rect 832 198 845 223
rect 1319 198 1332 244
rect 1378 238 1956 244
rect 1378 198 1391 238
rect 1943 198 1956 238
rect 2002 198 2083 244
rect 2605 220 4186 266
rect 5048 227 6857 289
rect 6953 273 6964 319
rect 7010 273 7163 319
rect 7209 273 7364 319
rect 7410 273 7603 319
rect 7649 273 7660 319
rect 518 166 662 177
rect 70 135 116 146
rect 294 139 340 152
rect 564 152 662 166
rect 928 152 1273 198
rect 2605 192 2651 220
rect 1437 152 1897 192
rect 2163 152 2536 192
rect 564 120 974 152
rect 518 106 974 120
rect 1227 146 2536 152
rect 2582 146 2651 192
rect 2760 163 2806 174
rect 1227 106 1483 146
rect 1851 106 2209 146
rect 294 60 340 93
rect 1020 95 1077 106
rect 0 49 1020 60
rect 1066 60 1077 95
rect 1631 60 1644 95
rect 1066 49 1644 60
rect 1690 60 1703 95
rect 2255 60 2268 95
rect 1690 49 2268 60
rect 2314 60 2327 95
rect 2760 60 2806 117
rect 2984 163 3030 220
rect 2984 106 3030 117
rect 3208 163 3254 174
rect 3208 60 3254 117
rect 3432 163 3478 220
rect 3432 106 3478 117
rect 3656 163 3702 174
rect 3656 60 3702 117
rect 3916 163 3962 220
rect 4351 219 7557 227
rect 3916 106 3962 117
rect 4140 163 4186 174
rect 4351 173 4364 219
rect 4410 173 4812 219
rect 4858 173 5260 219
rect 5306 173 5708 219
rect 5754 173 6156 219
rect 6202 173 6604 219
rect 6650 173 7052 219
rect 7098 173 7500 219
rect 7546 173 7557 219
rect 7724 192 7770 203
rect 4140 60 4186 117
rect 4577 81 4588 127
rect 4634 81 4645 127
rect 4577 60 4645 81
rect 5025 81 5036 127
rect 5082 81 5093 127
rect 5025 60 5093 81
rect 5473 81 5484 127
rect 5530 81 5541 127
rect 5473 60 5541 81
rect 5921 81 5932 127
rect 5978 81 5989 127
rect 5921 60 5989 81
rect 6369 81 6380 127
rect 6426 81 6437 127
rect 6369 60 6437 81
rect 6817 81 6828 127
rect 6874 81 6885 127
rect 6817 60 6885 81
rect 7265 81 7276 127
rect 7322 81 7333 127
rect 7265 60 7333 81
rect 7724 60 7770 146
rect 2314 49 7840 60
rect 0 -60 7840 49
<< labels >>
flabel metal1 s 0 724 7840 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 7724 174 7770 203 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 7500 601 7557 676 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 74 354 318 430 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 1026 354 1970 430 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 7045 601 7091 676 1 ZN
port 3 nsew default output
rlabel metal1 s 6595 601 6641 676 1 ZN
port 3 nsew default output
rlabel metal1 s 6151 601 6197 676 1 ZN
port 3 nsew default output
rlabel metal1 s 5702 601 5748 676 1 ZN
port 3 nsew default output
rlabel metal1 s 5251 601 5297 676 1 ZN
port 3 nsew default output
rlabel metal1 s 4805 601 4851 676 1 ZN
port 3 nsew default output
rlabel metal1 s 4364 601 4410 676 1 ZN
port 3 nsew default output
rlabel metal1 s 4364 485 7557 601 1 ZN
port 3 nsew default output
rlabel metal1 s 5790 289 5970 485 1 ZN
port 3 nsew default output
rlabel metal1 s 5048 227 6857 289 1 ZN
port 3 nsew default output
rlabel metal1 s 4351 173 7557 227 1 ZN
port 3 nsew default output
rlabel metal1 s 7704 689 7750 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7257 689 7325 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6810 689 6878 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6362 689 6430 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5914 689 5982 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5466 689 5534 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5016 689 5084 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4567 689 4635 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4136 689 4182 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3666 689 3712 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3199 689 3245 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2752 689 2798 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2270 689 2316 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1631 689 1703 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1009 689 1077 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 689 394 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7704 657 7750 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7257 657 7325 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6810 657 6878 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 6362 657 6430 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5914 657 5982 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5466 657 5534 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 5016 657 5084 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4567 657 4635 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4136 657 4182 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3666 657 3712 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3199 657 3245 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2752 657 2798 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2270 657 2316 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 326 657 394 689 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7704 540 7750 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 4136 540 4182 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3666 540 3712 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3199 540 3245 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2752 540 2798 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2270 540 2316 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7704 506 7750 540 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 7724 152 7770 174 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 152 4186 174 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3656 152 3702 174 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3208 152 3254 174 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2760 152 2806 174 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7724 127 7770 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 127 4186 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3656 127 3702 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3208 127 3254 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2760 127 2806 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 294 127 340 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7724 106 7770 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7265 106 7333 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6817 106 6885 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6369 106 6437 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5921 106 5989 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5473 106 5541 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5025 106 5093 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4577 106 4645 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 106 4186 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3656 106 3702 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3208 106 3254 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2760 106 2806 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 294 106 340 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7724 95 7770 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7265 95 7333 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6817 95 6885 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6369 95 6437 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5921 95 5989 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5473 95 5541 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5025 95 5093 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4577 95 4645 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 95 4186 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3656 95 3702 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3208 95 3254 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2760 95 2806 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1020 95 1077 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 294 95 340 106 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7724 60 7770 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 7265 60 7333 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6817 60 6885 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 6369 60 6437 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5921 60 5989 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5473 60 5541 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 5025 60 5093 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4577 60 4645 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 4140 60 4186 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3656 60 3702 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3208 60 3254 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2760 60 2806 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2255 60 2327 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1631 60 1703 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1020 60 1077 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 294 60 340 95 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 7840 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 7840 784
string GDS_END 569422
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 553772
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
