magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -50 448 50 453
rect -50 420 -45 448
rect -17 420 17 448
rect 45 420 50 448
rect -50 386 50 420
rect -50 358 -45 386
rect -17 358 17 386
rect 45 358 50 386
rect -50 324 50 358
rect -50 296 -45 324
rect -17 296 17 324
rect 45 296 50 324
rect -50 262 50 296
rect -50 234 -45 262
rect -17 234 17 262
rect 45 234 50 262
rect -50 200 50 234
rect -50 172 -45 200
rect -17 172 17 200
rect 45 172 50 200
rect -50 138 50 172
rect -50 110 -45 138
rect -17 110 17 138
rect 45 110 50 138
rect -50 76 50 110
rect -50 48 -45 76
rect -17 48 17 76
rect 45 48 50 76
rect -50 14 50 48
rect -50 -14 -45 14
rect -17 -14 17 14
rect 45 -14 50 14
rect -50 -48 50 -14
rect -50 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 50 -48
rect -50 -110 50 -76
rect -50 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 50 -110
rect -50 -172 50 -138
rect -50 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 50 -172
rect -50 -234 50 -200
rect -50 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 50 -234
rect -50 -296 50 -262
rect -50 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 50 -296
rect -50 -358 50 -324
rect -50 -386 -45 -358
rect -17 -386 17 -358
rect 45 -386 50 -358
rect -50 -420 50 -386
rect -50 -448 -45 -420
rect -17 -448 17 -420
rect 45 -448 50 -420
rect -50 -453 50 -448
<< via2 >>
rect -45 420 -17 448
rect 17 420 45 448
rect -45 358 -17 386
rect 17 358 45 386
rect -45 296 -17 324
rect 17 296 45 324
rect -45 234 -17 262
rect 17 234 45 262
rect -45 172 -17 200
rect 17 172 45 200
rect -45 110 -17 138
rect 17 110 45 138
rect -45 48 -17 76
rect 17 48 45 76
rect -45 -14 -17 14
rect 17 -14 45 14
rect -45 -76 -17 -48
rect 17 -76 45 -48
rect -45 -138 -17 -110
rect 17 -138 45 -110
rect -45 -200 -17 -172
rect 17 -200 45 -172
rect -45 -262 -17 -234
rect 17 -262 45 -234
rect -45 -324 -17 -296
rect 17 -324 45 -296
rect -45 -386 -17 -358
rect 17 -386 45 -358
rect -45 -448 -17 -420
rect 17 -448 45 -420
<< metal3 >>
rect -50 448 50 453
rect -50 420 -45 448
rect -17 420 17 448
rect 45 420 50 448
rect -50 386 50 420
rect -50 358 -45 386
rect -17 358 17 386
rect 45 358 50 386
rect -50 324 50 358
rect -50 296 -45 324
rect -17 296 17 324
rect 45 296 50 324
rect -50 262 50 296
rect -50 234 -45 262
rect -17 234 17 262
rect 45 234 50 262
rect -50 200 50 234
rect -50 172 -45 200
rect -17 172 17 200
rect 45 172 50 200
rect -50 138 50 172
rect -50 110 -45 138
rect -17 110 17 138
rect 45 110 50 138
rect -50 76 50 110
rect -50 48 -45 76
rect -17 48 17 76
rect 45 48 50 76
rect -50 14 50 48
rect -50 -14 -45 14
rect -17 -14 17 14
rect 45 -14 50 14
rect -50 -48 50 -14
rect -50 -76 -45 -48
rect -17 -76 17 -48
rect 45 -76 50 -48
rect -50 -110 50 -76
rect -50 -138 -45 -110
rect -17 -138 17 -110
rect 45 -138 50 -110
rect -50 -172 50 -138
rect -50 -200 -45 -172
rect -17 -200 17 -172
rect 45 -200 50 -172
rect -50 -234 50 -200
rect -50 -262 -45 -234
rect -17 -262 17 -234
rect 45 -262 50 -234
rect -50 -296 50 -262
rect -50 -324 -45 -296
rect -17 -324 17 -296
rect 45 -324 50 -296
rect -50 -358 50 -324
rect -50 -386 -45 -358
rect -17 -386 17 -358
rect 45 -386 50 -358
rect -50 -420 50 -386
rect -50 -448 -45 -420
rect -17 -448 17 -420
rect 45 -448 50 -420
rect -50 -453 50 -448
<< properties >>
string GDS_END 1104394
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1102342
<< end >>
