magic
tech gf180mcuC
timestamp 1666464484
<< properties >>
string GDS_END 14432458
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 14323910
<< end >>
