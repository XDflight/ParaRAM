magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 341 89 414
rect 193 341 313 414
use pmos_5p04310589983266_64x8m81  pmos_5p04310589983266_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 552 462
<< properties >>
string GDS_END 214494
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 214116
<< end >>
