magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -60 -407 1259 1742
<< pmos >>
rect 206 507 994 1606
<< pdiff >>
rect 81 1563 206 1606
rect 81 1517 127 1563
rect 173 1517 206 1563
rect 81 1402 206 1517
rect 81 1356 127 1402
rect 173 1356 206 1402
rect 81 1242 206 1356
rect 81 1196 127 1242
rect 173 1196 206 1242
rect 81 1082 206 1196
rect 81 1036 127 1082
rect 173 1036 206 1082
rect 81 921 206 1036
rect 81 875 127 921
rect 173 875 206 921
rect 81 759 206 875
rect 81 713 127 759
rect 173 713 206 759
rect 81 596 206 713
rect 81 550 127 596
rect 173 550 206 596
rect 81 507 206 550
rect 994 1563 1119 1606
rect 994 1517 1027 1563
rect 1073 1517 1119 1563
rect 994 1402 1119 1517
rect 994 1356 1027 1402
rect 1073 1356 1119 1402
rect 994 1242 1119 1356
rect 994 1196 1027 1242
rect 1073 1196 1119 1242
rect 994 1082 1119 1196
rect 994 1036 1027 1082
rect 1073 1036 1119 1082
rect 994 921 1119 1036
rect 994 875 1027 921
rect 1073 875 1119 921
rect 994 759 1119 875
rect 994 713 1027 759
rect 1073 713 1119 759
rect 994 596 1119 713
rect 994 550 1027 596
rect 1073 550 1119 596
rect 994 507 1119 550
<< pdiffc >>
rect 127 1517 173 1563
rect 127 1356 173 1402
rect 127 1196 173 1242
rect 127 1036 173 1082
rect 127 875 173 921
rect 127 713 173 759
rect 127 550 173 596
rect 1027 1517 1073 1563
rect 1027 1356 1073 1402
rect 1027 1196 1073 1242
rect 1027 1036 1073 1082
rect 1027 875 1073 921
rect 1027 713 1073 759
rect 1027 550 1073 596
<< psubdiff >>
rect 49 2070 1150 2124
rect 49 2024 255 2070
rect 301 2024 419 2070
rect 465 2024 582 2070
rect 628 2024 745 2070
rect 791 2024 909 2070
rect 955 2024 1150 2070
rect 49 1969 1150 2024
<< nsubdiff >>
rect 83 243 1116 297
rect 83 197 255 243
rect 301 197 419 243
rect 465 197 582 243
rect 628 197 745 243
rect 791 197 909 243
rect 955 197 1116 243
rect 83 78 1116 197
<< psubdiffcont >>
rect 255 2024 301 2070
rect 419 2024 465 2070
rect 582 2024 628 2070
rect 745 2024 791 2070
rect 909 2024 955 2070
<< nsubdiffcont >>
rect 255 197 301 243
rect 419 197 465 243
rect 582 197 628 243
rect 745 197 791 243
rect 909 197 955 243
<< polysilicon >>
rect 206 1764 994 1808
rect 206 1718 333 1764
rect 379 1718 496 1764
rect 542 1718 660 1764
rect 706 1718 823 1764
rect 869 1718 994 1764
rect 206 1606 994 1718
rect 206 436 994 507
<< polycontact >>
rect 333 1718 379 1764
rect 496 1718 542 1764
rect 660 1718 706 1764
rect 823 1718 869 1764
<< metal1 >>
rect 49 2070 1150 2124
rect 49 2035 255 2070
rect 49 1983 124 2035
rect 176 2024 255 2035
rect 301 2024 419 2070
rect 465 2024 582 2070
rect 628 2024 745 2070
rect 791 2024 909 2070
rect 955 2024 1150 2070
rect 176 1983 1150 2024
rect 49 1824 1150 1983
rect 49 1772 124 1824
rect 176 1772 1150 1824
rect 49 1764 1150 1772
rect 49 1718 333 1764
rect 379 1718 496 1764
rect 542 1718 660 1764
rect 706 1718 823 1764
rect 869 1718 1150 1764
rect 49 1684 1150 1718
rect 83 1563 216 1597
rect 83 1517 127 1563
rect 173 1517 216 1563
rect 83 1402 216 1517
rect 83 1356 127 1402
rect 173 1356 216 1402
rect 83 1336 216 1356
rect 983 1563 1116 1597
rect 983 1517 1027 1563
rect 1073 1517 1116 1563
rect 983 1402 1116 1517
rect 983 1356 1027 1402
rect 1073 1356 1116 1402
rect 983 1336 1116 1356
rect 83 1298 217 1336
rect 83 1246 124 1298
rect 176 1246 217 1298
rect 83 1242 217 1246
rect 83 1196 127 1242
rect 173 1196 217 1242
rect 83 1087 217 1196
rect 83 1035 124 1087
rect 176 1035 217 1087
rect 83 921 217 1035
rect 83 875 127 921
rect 173 875 217 921
rect 83 823 124 875
rect 176 823 217 875
rect 83 759 217 823
rect 83 713 127 759
rect 173 713 217 759
rect 83 664 217 713
rect 83 612 124 664
rect 176 612 217 664
rect 83 596 217 612
rect 83 550 127 596
rect 173 574 217 596
rect 983 1298 1117 1336
rect 983 1246 1024 1298
rect 1076 1246 1117 1298
rect 983 1242 1117 1246
rect 983 1196 1027 1242
rect 1073 1196 1117 1242
rect 983 1087 1117 1196
rect 983 1035 1024 1087
rect 1076 1035 1117 1087
rect 983 921 1117 1035
rect 983 875 1027 921
rect 1073 875 1117 921
rect 983 823 1024 875
rect 1076 823 1117 875
rect 983 759 1117 823
rect 983 713 1027 759
rect 1073 713 1117 759
rect 983 664 1117 713
rect 983 612 1024 664
rect 1076 612 1117 664
rect 983 596 1117 612
rect 173 550 216 574
rect 83 515 216 550
rect 983 550 1027 596
rect 1073 574 1117 596
rect 1073 550 1116 574
rect 983 515 1116 550
rect 83 243 1116 297
rect 83 197 255 243
rect 301 197 419 243
rect 465 197 582 243
rect 628 197 745 243
rect 791 197 909 243
rect 955 197 1116 243
rect 83 78 1116 197
<< via1 >>
rect 124 1983 176 2035
rect 124 1772 176 1824
rect 124 1246 176 1298
rect 124 1082 176 1087
rect 124 1036 127 1082
rect 127 1036 173 1082
rect 173 1036 176 1082
rect 124 1035 176 1036
rect 124 823 176 875
rect 124 612 176 664
rect 1024 1246 1076 1298
rect 1024 1082 1076 1087
rect 1024 1036 1027 1082
rect 1027 1036 1073 1082
rect 1073 1036 1076 1082
rect 1024 1035 1076 1036
rect 1024 823 1076 875
rect 1024 612 1076 664
<< metal2 >>
rect 83 2037 217 2074
rect 83 1981 122 2037
rect 178 1981 217 2037
rect 83 1826 217 1981
rect 83 1770 122 1826
rect 178 1770 217 1826
rect 83 1734 217 1770
rect 49 1300 1150 1395
rect 49 1298 1022 1300
rect 49 1246 124 1298
rect 176 1246 1022 1298
rect 49 1244 1022 1246
rect 1078 1244 1150 1300
rect 49 1089 1150 1244
rect 49 1087 1022 1089
rect 49 1035 124 1087
rect 176 1035 1022 1087
rect 49 1033 1022 1035
rect 1078 1033 1150 1089
rect 49 877 1150 1033
rect 49 875 1022 877
rect 49 823 124 875
rect 176 823 1022 875
rect 49 821 1022 823
rect 1078 821 1150 877
rect 49 666 1150 821
rect 49 664 1022 666
rect 49 612 124 664
rect 176 612 1022 664
rect 49 610 1022 612
rect 1078 610 1150 666
rect 49 515 1150 610
<< via2 >>
rect 122 2035 178 2037
rect 122 1983 124 2035
rect 124 1983 176 2035
rect 176 1983 178 2035
rect 122 1981 178 1983
rect 122 1824 178 1826
rect 122 1772 124 1824
rect 124 1772 176 1824
rect 176 1772 178 1824
rect 122 1770 178 1772
rect 1022 1298 1078 1300
rect 1022 1246 1024 1298
rect 1024 1246 1076 1298
rect 1076 1246 1078 1298
rect 1022 1244 1078 1246
rect 1022 1087 1078 1089
rect 1022 1035 1024 1087
rect 1024 1035 1076 1087
rect 1076 1035 1078 1087
rect 1022 1033 1078 1035
rect 1022 875 1078 877
rect 1022 823 1024 875
rect 1024 823 1076 875
rect 1076 823 1078 875
rect 1022 821 1078 823
rect 1022 664 1078 666
rect 1022 612 1024 664
rect 1024 612 1076 664
rect 1076 612 1078 664
rect 1022 610 1078 612
<< metal3 >>
rect 49 2037 250 3251
rect 49 1981 122 2037
rect 178 1981 250 2037
rect 49 1826 250 1981
rect 49 1770 122 1826
rect 178 1770 250 1826
rect 49 -1 250 1770
rect 509 -1 711 2203
rect 949 1300 1150 2204
rect 949 1244 1022 1300
rect 1078 1244 1150 1300
rect 949 1089 1150 1244
rect 949 1033 1022 1089
rect 1078 1033 1150 1089
rect 949 877 1150 1033
rect 949 821 1022 877
rect 1078 821 1150 877
rect 949 666 1150 821
rect 949 610 1022 666
rect 1078 610 1150 666
rect 949 -1 1150 610
use M1_NACTIVE$$2042_R270_64x8m81  M1_NACTIVE$$2042_R270_64x8m81_0
timestamp 1666464484
transform 1 0 605 0 1 220
box 0 0 1 1
use M1_PACTIVE$$2042_R270_64x8m81  M1_PACTIVE$$2042_R270_64x8m81_0
timestamp 1666464484
transform 1 0 605 0 1 2047
box 0 0 1 1
use M1_POLY2$$2043_R270_64x8m81  M1_POLY2$$2043_R270_64x8m81_0
timestamp 1666464484
transform 1 0 601 0 1 1741
box 0 0 1 1
use M2_M1$$204396588_R270_64x8m81  M2_M1$$204396588_R270_64x8m81_0
timestamp 1666464484
transform 1 0 150 0 1 955
box 0 0 1 1
use M2_M1$$204396588_R270_64x8m81  M2_M1$$204396588_R270_64x8m81_1
timestamp 1666464484
transform 1 0 1050 0 1 955
box 0 0 1 1
use M3_M2$$204397612_R270_64x8m81  M3_M2$$204397612_R270_64x8m81_0
timestamp 1666464484
transform 1 0 1050 0 1 955
box 0 0 1 1
<< properties >>
string GDS_END 1331620
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1328862
<< end >>
