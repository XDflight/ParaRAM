magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 1878 870
<< pwell >>
rect -86 -86 1878 352
<< mvnmos >>
rect 124 68 324 232
rect 572 68 772 232
rect 1020 68 1220 232
rect 1468 68 1668 232
<< mvpmos >>
rect 124 472 324 716
rect 572 472 772 716
rect 1020 472 1220 716
rect 1468 472 1668 716
<< mvndiff >>
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 324 192 412 232
rect 324 146 353 192
rect 399 146 412 192
rect 324 68 412 146
rect 484 192 572 232
rect 484 146 497 192
rect 543 146 572 192
rect 484 68 572 146
rect 772 192 860 232
rect 772 146 801 192
rect 847 146 860 192
rect 772 68 860 146
rect 932 192 1020 232
rect 932 146 945 192
rect 991 146 1020 192
rect 932 68 1020 146
rect 1220 192 1308 232
rect 1220 146 1249 192
rect 1295 146 1308 192
rect 1220 68 1308 146
rect 1380 192 1468 232
rect 1380 146 1393 192
rect 1439 146 1468 192
rect 1380 68 1468 146
rect 1668 192 1756 232
rect 1668 146 1697 192
rect 1743 146 1756 192
rect 1668 68 1756 146
<< mvpdiff >>
rect 36 657 124 716
rect 36 517 49 657
rect 95 517 124 657
rect 36 472 124 517
rect 324 657 412 716
rect 324 517 353 657
rect 399 517 412 657
rect 324 472 412 517
rect 484 657 572 716
rect 484 517 497 657
rect 543 517 572 657
rect 484 472 572 517
rect 772 657 860 716
rect 772 517 801 657
rect 847 517 860 657
rect 772 472 860 517
rect 932 657 1020 716
rect 932 517 945 657
rect 991 517 1020 657
rect 932 472 1020 517
rect 1220 657 1308 716
rect 1220 517 1249 657
rect 1295 517 1308 657
rect 1220 472 1308 517
rect 1380 657 1468 716
rect 1380 517 1393 657
rect 1439 517 1468 657
rect 1380 472 1468 517
rect 1668 657 1756 716
rect 1668 517 1697 657
rect 1743 517 1756 657
rect 1668 472 1756 517
<< mvndiffc >>
rect 49 146 95 192
rect 353 146 399 192
rect 497 146 543 192
rect 801 146 847 192
rect 945 146 991 192
rect 1249 146 1295 192
rect 1393 146 1439 192
rect 1697 146 1743 192
<< mvpdiffc >>
rect 49 517 95 657
rect 353 517 399 657
rect 497 517 543 657
rect 801 517 847 657
rect 945 517 991 657
rect 1249 517 1295 657
rect 1393 517 1439 657
rect 1697 517 1743 657
<< polysilicon >>
rect 124 716 324 760
rect 572 716 772 760
rect 1020 716 1220 760
rect 1468 716 1668 760
rect 124 438 324 472
rect 124 392 160 438
rect 300 392 324 438
rect 124 375 324 392
rect 572 438 772 472
rect 572 392 608 438
rect 748 392 772 438
rect 572 375 772 392
rect 1020 438 1220 472
rect 1020 392 1056 438
rect 1196 392 1220 438
rect 1020 375 1220 392
rect 1468 438 1668 472
rect 1468 392 1504 438
rect 1644 392 1668 438
rect 1468 375 1668 392
rect 124 311 324 324
rect 124 265 152 311
rect 292 265 324 311
rect 124 232 324 265
rect 572 311 772 324
rect 572 265 600 311
rect 740 265 772 311
rect 572 232 772 265
rect 1020 311 1220 324
rect 1020 265 1048 311
rect 1188 265 1220 311
rect 1020 232 1220 265
rect 1468 311 1668 324
rect 1468 265 1496 311
rect 1636 265 1668 311
rect 1468 232 1668 265
rect 124 24 324 68
rect 572 24 772 68
rect 1020 24 1220 68
rect 1468 24 1668 68
<< polycontact >>
rect 160 392 300 438
rect 608 392 748 438
rect 1056 392 1196 438
rect 1504 392 1644 438
rect 152 265 292 311
rect 600 265 740 311
rect 1048 265 1188 311
rect 1496 265 1636 311
<< metal1 >>
rect 0 724 1792 844
rect 49 657 95 678
rect 49 311 95 517
rect 353 657 399 724
rect 353 498 399 517
rect 497 657 543 678
rect 146 392 160 438
rect 300 392 399 438
rect 49 265 152 311
rect 292 265 304 311
rect 49 192 95 214
rect 49 60 95 146
rect 353 192 399 392
rect 497 311 543 517
rect 801 657 847 724
rect 801 498 847 517
rect 945 657 991 678
rect 594 392 608 438
rect 748 392 847 438
rect 497 265 600 311
rect 740 265 752 311
rect 353 106 399 146
rect 497 192 543 214
rect 497 60 543 146
rect 801 192 847 392
rect 945 311 991 517
rect 1249 657 1295 724
rect 1249 498 1295 517
rect 1393 657 1439 678
rect 1042 392 1056 438
rect 1196 392 1295 438
rect 945 265 1048 311
rect 1188 265 1200 311
rect 801 106 847 146
rect 945 192 991 214
rect 945 60 991 146
rect 1249 192 1295 392
rect 1393 311 1439 517
rect 1697 657 1743 724
rect 1697 498 1743 517
rect 1490 392 1504 438
rect 1644 392 1743 438
rect 1393 265 1496 311
rect 1636 265 1648 311
rect 1249 106 1295 146
rect 1393 192 1439 214
rect 1393 60 1439 146
rect 1697 192 1743 392
rect 1697 106 1743 146
rect 0 -60 1792 60
<< labels >>
flabel metal1 s 0 724 1792 844 0 FreeSans 400 0 0 0 VDD
port 1 nsew power bidirectional abutment
flabel metal1 s 1393 60 1439 214 0 FreeSans 400 0 0 0 VSS
port 4 nsew ground bidirectional abutment
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 1697 498 1743 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 498 1295 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 498 847 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 1 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 945 60 991 214 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 214 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 214 1 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1792 60 1 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 784
string GDS_END 1143332
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1137820
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
