magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 191 88 264
rect -31 -73 88 -1
use nmos_5p0431059054878_128x8m81  nmos_5p0431059054878_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 208 236
<< properties >>
string GDS_END 232130
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 231880
<< end >>
