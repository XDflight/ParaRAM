magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
use 018SRAM_cell1_64x8m81  018SRAM_cell1_64x8m81_0
timestamp 1666464484
transform 1 0 0 0 -1 450
box -34 -34 334 484
use 018SRAM_cell1_64x8m81  018SRAM_cell1_64x8m81_1
timestamp 1666464484
transform 1 0 0 0 1 450
box -34 -34 334 484
<< properties >>
string GDS_END 567592
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 567490
<< end >>
