magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 1206 870
<< pwell >>
rect -86 -86 1206 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 796 68 916 232
<< mvpmos >>
rect 144 472 244 716
rect 348 472 448 716
rect 592 519 692 716
rect 796 519 896 716
<< mvndiff >>
rect 36 167 124 232
rect 36 121 49 167
rect 95 121 124 167
rect 36 68 124 121
rect 244 167 348 232
rect 244 121 273 167
rect 319 121 348 167
rect 244 68 348 121
rect 468 167 572 232
rect 468 121 497 167
rect 543 121 572 167
rect 468 68 572 121
rect 692 68 796 232
rect 916 167 1004 232
rect 916 121 945 167
rect 991 121 1004 167
rect 916 68 1004 121
<< mvpdiff >>
rect 46 641 144 716
rect 46 595 59 641
rect 105 595 144 641
rect 46 472 144 595
rect 244 472 348 716
rect 448 586 592 716
rect 448 540 497 586
rect 543 540 592 586
rect 448 519 592 540
rect 692 703 796 716
rect 692 657 721 703
rect 767 657 796 703
rect 692 519 796 657
rect 896 586 986 716
rect 896 540 927 586
rect 973 540 986 586
rect 896 519 986 540
rect 448 472 528 519
<< mvndiffc >>
rect 49 121 95 167
rect 273 121 319 167
rect 497 121 543 167
rect 945 121 991 167
<< mvpdiffc >>
rect 59 595 105 641
rect 497 540 543 586
rect 721 657 767 703
rect 927 540 973 586
<< polysilicon >>
rect 144 716 244 760
rect 348 716 448 760
rect 592 716 692 760
rect 796 716 896 760
rect 144 402 244 472
rect 124 368 244 402
rect 124 322 147 368
rect 193 322 244 368
rect 124 232 244 322
rect 348 402 448 472
rect 592 415 692 519
rect 592 402 611 415
rect 348 368 468 402
rect 348 322 371 368
rect 417 322 468 368
rect 348 232 468 322
rect 572 369 611 402
rect 657 369 692 415
rect 572 232 692 369
rect 796 415 896 519
rect 796 369 823 415
rect 869 402 896 415
rect 869 369 916 402
rect 796 232 916 369
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 796 24 916 68
<< polycontact >>
rect 147 322 193 368
rect 371 322 417 368
rect 611 369 657 415
rect 823 369 869 415
<< metal1 >>
rect 0 724 1120 844
rect 59 641 105 724
rect 710 703 778 724
rect 59 584 105 595
rect 151 632 658 678
rect 710 657 721 703
rect 767 657 778 703
rect 151 538 197 632
rect 612 611 658 632
rect 824 632 1090 678
rect 824 611 870 632
rect 486 540 497 586
rect 543 540 554 586
rect 612 565 870 611
rect 49 492 197 538
rect 248 519 554 540
rect 916 540 927 586
rect 973 540 984 586
rect 916 519 984 540
rect 49 167 95 492
rect 248 473 984 519
rect 49 110 95 121
rect 141 368 200 446
rect 141 322 147 368
rect 193 322 200 368
rect 141 110 200 322
rect 248 167 319 473
rect 248 121 273 167
rect 248 110 319 121
rect 365 368 424 427
rect 365 322 371 368
rect 417 322 424 368
rect 365 110 424 322
rect 472 415 674 424
rect 472 369 611 415
rect 657 369 674 415
rect 472 360 674 369
rect 730 415 994 424
rect 730 369 823 415
rect 869 369 994 415
rect 730 360 994 369
rect 472 232 532 360
rect 730 312 788 360
rect 578 248 788 312
rect 1044 274 1090 632
rect 848 228 1090 274
rect 848 167 894 228
rect 486 121 497 167
rect 543 121 894 167
rect 848 120 894 121
rect 945 167 991 178
rect 945 60 991 121
rect 0 -60 1120 60
<< labels >>
flabel metal1 s 472 360 674 424 0 FreeSans 400 0 0 0 B
port 3 nsew default input
flabel metal1 s 730 360 994 424 0 FreeSans 400 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 724 1120 844 0 FreeSans 400 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 945 60 991 178 0 FreeSans 400 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 916 540 984 586 0 FreeSans 400 0 0 0 ZN
port 5 nsew default output
flabel metal1 s 365 110 424 427 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 141 110 200 446 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 472 232 532 360 1 B
port 3 nsew default input
rlabel metal1 s 730 312 788 360 1 C
port 4 nsew default input
rlabel metal1 s 578 248 788 312 1 C
port 4 nsew default input
rlabel metal1 s 486 540 554 586 1 ZN
port 5 nsew default output
rlabel metal1 s 916 519 984 540 1 ZN
port 5 nsew default output
rlabel metal1 s 248 519 554 540 1 ZN
port 5 nsew default output
rlabel metal1 s 248 473 984 519 1 ZN
port 5 nsew default output
rlabel metal1 s 248 110 319 473 1 ZN
port 5 nsew default output
rlabel metal1 s 710 657 778 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 657 105 724 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 59 584 105 657 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -60 1120 60 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 784
string GDS_END 90518
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 87160
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
