magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect 27097 35977 28629 96310
rect 55930 35977 57389 96310
rect 85432 578 85816 96702
<< metal1 >>
rect 0 403 1000 96694
<< metal2 >>
rect 424 403 1424 96149
<< metal3 >>
rect 424 0 1424 2232
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_0
timestamp 1666464484
transform -1 0 85672 0 1 96288
box -42 -42 85602 414
use M1_PSUB4310591302043_512x8m81  M1_PSUB4310591302043_512x8m81_1
timestamp 1666464484
transform -1 0 85672 0 1 620
box -42 -42 85602 414
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_0
timestamp 1666464484
transform 1 0 85474 0 1 1140
box -42 -42 342 95042
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_1
timestamp 1666464484
transform 1 0 27139 0 1 1140
box -42 -42 342 95042
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_2
timestamp 1666464484
transform 1 0 57047 0 1 1140
box -42 -42 342 95042
use M1_PSUB4310591302044_512x8m81  M1_PSUB4310591302044_512x8m81_3
timestamp 1666464484
transform 1 0 112 0 1 1140
box -42 -42 342 95042
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_0
timestamp 1666464484
transform 1 0 56123 0 1 36019
box -42 -42 842 60142
use M1_PSUB4310591302045_512x8m81  M1_PSUB4310591302045_512x8m81_1
timestamp 1666464484
transform 1 0 27563 0 1 36019
box -42 -42 842 60142
use M1_PSUB4310591302046_512x8m81  M1_PSUB4310591302046_512x8m81_0
timestamp 1666464484
transform 1 0 27563 0 1 34197
box -42 -42 29342 442
<< labels >>
flabel metal3 s 924 178 924 178 0 FreeSans 2000 0 0 0 VDD
port 1 nsew
<< properties >>
string GDS_END 2641600
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2640290
string path 4.620 11.160 4.620 0.000 
<< end >>
