magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -19 247 19 253
rect -19 -247 -13 247
rect 13 -247 19 247
rect -19 -253 19 -247
<< via1 >>
rect -13 -247 13 247
<< metal2 >>
rect -19 247 19 253
rect -19 -247 -13 247
rect 13 -247 19 247
rect -19 -253 19 -247
<< properties >>
string GDS_END 514354
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 513582
<< end >>
