magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 4256 844
rect 252 569 320 724
rect 1050 636 1118 724
rect 1514 670 1582 724
rect 141 119 206 430
rect 273 60 319 228
rect 365 119 430 430
rect 682 359 1017 443
rect 1093 359 1326 440
rect 1059 60 1127 215
rect 1556 60 1602 209
rect 2586 599 2654 724
rect 2596 60 2664 217
rect 3450 569 3518 724
rect 3947 492 3993 724
rect 3525 60 3571 136
rect 3937 60 3983 199
rect 4158 123 4230 673
rect 0 -60 4256 60
<< obsm1 >>
rect 49 523 95 603
rect 1175 624 1464 664
rect 1674 624 2003 670
rect 1175 618 1720 624
rect 1175 587 1221 618
rect 606 541 1221 587
rect 1418 578 1720 618
rect 1317 532 1363 572
rect 49 477 555 523
rect 1317 486 1720 532
rect 49 158 95 477
rect 509 325 555 477
rect 885 261 1264 307
rect 885 215 931 261
rect 654 169 931 215
rect 1218 152 1264 261
rect 1372 255 1418 486
rect 1674 375 1720 486
rect 1780 410 1826 572
rect 1957 538 2003 624
rect 2065 630 2498 678
rect 2065 410 2111 630
rect 1780 364 2111 410
rect 1350 198 1418 255
rect 1464 261 1721 307
rect 1464 152 1510 261
rect 1218 106 1510 152
rect 1675 152 1721 261
rect 1813 255 1859 364
rect 2171 340 2217 574
rect 2452 553 2498 630
rect 2734 632 3249 678
rect 2734 553 2780 632
rect 2452 506 2780 553
rect 2865 460 2911 574
rect 2440 414 2911 460
rect 2171 294 2793 340
rect 1813 198 1881 255
rect 1968 152 2014 228
rect 2192 160 2238 294
rect 1675 106 2014 152
rect 2865 160 2911 414
rect 2957 252 3003 632
rect 3089 355 3135 574
rect 3181 414 3249 632
rect 3301 463 3634 510
rect 3301 355 3347 463
rect 3089 308 3347 355
rect 3566 334 3634 463
rect 3693 402 3739 590
rect 3693 356 4108 402
rect 3089 160 3135 308
rect 3393 246 3439 320
rect 3793 246 3839 356
rect 3393 199 3839 246
rect 3793 152 3839 199
<< labels >>
rlabel metal1 s 682 359 1017 443 6 D
port 1 nsew default input
rlabel metal1 s 141 119 206 430 6 SE
port 2 nsew default input
rlabel metal1 s 365 119 430 430 6 SI
port 3 nsew default input
rlabel metal1 s 1093 359 1326 440 6 CLK
port 4 nsew clock input
rlabel metal1 s 4158 123 4230 673 6 Q
port 5 nsew default output
rlabel metal1 s 0 724 4256 844 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 670 3993 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 670 3518 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 670 2654 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1514 670 1582 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 670 1118 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 724 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 636 3993 670 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 636 3518 670 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 636 2654 670 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1050 636 1118 670 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 636 320 670 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 599 3993 636 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 599 3518 636 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2586 599 2654 636 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 599 320 636 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 569 3993 599 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3450 569 3518 599 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 599 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3947 492 3993 569 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 217 319 228 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 215 2664 217 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 215 319 217 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 209 2664 215 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 209 1127 215 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 209 319 215 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 199 2664 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 199 1602 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 199 1127 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 199 319 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3937 136 3983 199 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 136 2664 199 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 136 1602 199 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 136 1127 199 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 136 319 199 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3937 60 3983 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3525 60 3571 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2596 60 2664 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1556 60 1602 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1059 60 1127 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 136 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4256 60 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4256 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 186850
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 178018
<< end >>
