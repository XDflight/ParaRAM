magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 3472 844
rect 262 586 330 724
rect 661 637 707 724
rect 130 354 318 430
rect 262 60 330 210
rect 630 60 698 218
rect 914 242 995 542
rect 1526 540 1594 724
rect 2525 527 2571 724
rect 2873 527 2919 724
rect 3066 466 3282 595
rect 3333 527 3379 724
rect 1558 60 1626 117
rect 2497 60 2543 221
rect 3206 204 3282 466
rect 2885 60 2931 178
rect 3090 110 3282 204
rect 3333 60 3379 194
rect 0 -60 3472 60
<< obsm1 >>
rect 69 540 115 631
rect 383 596 615 643
rect 383 540 429 596
rect 569 577 615 596
rect 778 632 1318 678
rect 778 577 824 632
rect 69 494 429 540
rect 383 302 429 494
rect 477 465 523 542
rect 569 530 824 577
rect 477 418 815 465
rect 769 311 815 418
rect 49 256 429 302
rect 497 265 815 311
rect 49 162 95 256
rect 497 162 543 265
rect 769 152 815 265
rect 1122 494 1190 586
rect 1728 632 2266 678
rect 1065 448 1682 494
rect 1065 198 1134 448
rect 1728 402 1774 632
rect 1233 356 1774 402
rect 1233 152 1279 356
rect 1825 310 1894 586
rect 1426 264 1894 310
rect 1826 172 1894 264
rect 1944 245 1990 632
rect 2050 426 2118 586
rect 2050 379 2670 426
rect 2050 172 2118 379
rect 2729 368 2775 606
rect 2729 326 3113 368
rect 2354 300 3113 326
rect 2354 280 2774 300
rect 769 106 1279 152
rect 2721 161 2774 280
<< labels >>
rlabel metal1 s 914 242 995 542 6 D
port 1 nsew default input
rlabel metal1 s 130 354 318 430 6 CLK
port 2 nsew clock input
rlabel metal1 s 3066 466 3282 595 6 Q
port 3 nsew default output
rlabel metal1 s 3206 204 3282 466 6 Q
port 3 nsew default output
rlabel metal1 s 3090 110 3282 204 6 Q
port 3 nsew default output
rlabel metal1 s 0 724 3472 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 637 3379 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 637 2919 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 637 2571 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 637 1594 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 661 637 707 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 262 637 330 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 586 3379 637 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 586 2919 637 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 586 2571 637 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 586 1594 637 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 262 586 330 637 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 540 3379 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 540 2919 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 540 2571 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1526 540 1594 586 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3333 527 3379 540 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2873 527 2919 540 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2525 527 2571 540 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2497 218 2543 221 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2497 210 2543 218 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 630 210 698 218 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2497 194 2543 210 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 630 194 698 210 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 194 330 210 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3333 178 3379 194 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2497 178 2543 194 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 630 178 698 194 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 178 330 194 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3333 117 3379 178 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2885 117 2931 178 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2497 117 2543 178 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 630 117 698 178 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 117 330 178 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3333 60 3379 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2885 60 2931 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2497 60 2543 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1558 60 1626 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 630 60 698 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 117 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3472 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3472 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 963166
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 955882
<< end >>
