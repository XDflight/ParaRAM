magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -81 292 81 298
rect -81 266 -75 292
rect -49 266 -13 292
rect 13 266 49 292
rect 75 266 81 292
rect -81 230 81 266
rect -81 204 -75 230
rect -49 204 -13 230
rect 13 204 49 230
rect 75 204 81 230
rect -81 168 81 204
rect -81 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 81 168
rect -81 106 81 142
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -142 81 -106
rect -81 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 81 -142
rect -81 -204 81 -168
rect -81 -230 -75 -204
rect -49 -230 -13 -204
rect 13 -230 49 -204
rect 75 -230 81 -204
rect -81 -266 81 -230
rect -81 -292 -75 -266
rect -49 -292 -13 -266
rect 13 -292 49 -266
rect 75 -292 81 -266
rect -81 -298 81 -292
<< via1 >>
rect -75 266 -49 292
rect -13 266 13 292
rect 49 266 75 292
rect -75 204 -49 230
rect -13 204 13 230
rect 49 204 75 230
rect -75 142 -49 168
rect -13 142 13 168
rect 49 142 75 168
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
rect -75 -168 -49 -142
rect -13 -168 13 -142
rect 49 -168 75 -142
rect -75 -230 -49 -204
rect -13 -230 13 -204
rect 49 -230 75 -204
rect -75 -292 -49 -266
rect -13 -292 13 -266
rect 49 -292 75 -266
<< metal2 >>
rect -81 292 81 298
rect -81 266 -75 292
rect -49 266 -13 292
rect 13 266 49 292
rect 75 266 81 292
rect -81 230 81 266
rect -81 204 -75 230
rect -49 204 -13 230
rect 13 204 49 230
rect 75 204 81 230
rect -81 168 81 204
rect -81 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 81 168
rect -81 106 81 142
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -142 81 -106
rect -81 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 81 -142
rect -81 -204 81 -168
rect -81 -230 -75 -204
rect -49 -230 -13 -204
rect 13 -230 49 -204
rect 75 -230 81 -204
rect -81 -266 81 -230
rect -81 -292 -75 -266
rect -49 -292 -13 -266
rect 13 -292 49 -266
rect 75 -292 81 -266
rect -81 -298 81 -292
<< properties >>
string GDS_END 728960
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 726908
<< end >>
