magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect 495 6267 719 7462
rect 495 6211 516 6267
rect 572 6211 640 6267
rect 696 6211 719 6267
rect 495 6143 719 6211
rect 495 6087 516 6143
rect 572 6087 640 6143
rect 696 6087 719 6143
rect 495 6019 719 6087
rect 495 5963 516 6019
rect 572 5963 640 6019
rect 696 5963 719 6019
rect -8 4667 216 5604
rect -8 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 216 4667
rect -8 4543 216 4611
rect -8 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 216 4543
rect -8 4419 216 4487
rect -8 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 216 4419
rect -8 2115 216 4363
rect 495 3065 719 5963
rect 1011 4667 1235 5605
rect 1011 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1235 4667
rect 1011 4543 1235 4611
rect 1011 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1235 4543
rect 1011 4419 1235 4487
rect 1011 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1235 4419
rect 1011 2115 1235 4363
<< via2 >>
rect 516 6211 572 6267
rect 640 6211 696 6267
rect 516 6087 572 6143
rect 640 6087 696 6143
rect 516 5963 572 6019
rect 640 5963 696 6019
rect 16 4611 72 4667
rect 140 4611 196 4667
rect 16 4487 72 4543
rect 140 4487 196 4543
rect 16 4363 72 4419
rect 140 4363 196 4419
rect 1033 4611 1089 4667
rect 1157 4611 1213 4667
rect 1033 4487 1089 4543
rect 1157 4487 1213 4543
rect 1033 4363 1089 4419
rect 1157 4363 1213 4419
<< metal3 >>
rect 506 6267 706 6277
rect 506 6211 516 6267
rect 572 6211 640 6267
rect 696 6211 706 6267
rect 506 6143 706 6211
rect 506 6087 516 6143
rect 572 6087 640 6143
rect 696 6087 706 6143
rect 506 6019 706 6087
rect 506 5963 516 6019
rect 572 5963 640 6019
rect 696 5963 706 6019
rect 506 5953 706 5963
rect 6 4667 206 4677
rect 6 4611 16 4667
rect 72 4611 140 4667
rect 196 4611 206 4667
rect 6 4543 206 4611
rect 6 4487 16 4543
rect 72 4487 140 4543
rect 196 4487 206 4543
rect 6 4419 206 4487
rect 6 4363 16 4419
rect 72 4363 140 4419
rect 196 4363 206 4419
rect 6 4353 206 4363
rect 1023 4667 1223 4677
rect 1023 4611 1033 4667
rect 1089 4611 1157 4667
rect 1213 4611 1223 4667
rect 1023 4543 1223 4611
rect 1023 4487 1033 4543
rect 1089 4487 1157 4543
rect 1213 4487 1223 4543
rect 1023 4419 1223 4487
rect 1023 4363 1033 4419
rect 1089 4363 1157 4419
rect 1213 4363 1223 4419
rect 1023 4353 1223 4363
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_0
timestamp 1666464484
transform 1 0 1120 0 1 2602
box -100 -472 100 472
use M2_M14310590878176_256x8m81  M2_M14310590878176_256x8m81_1
timestamp 1666464484
transform 1 0 103 0 1 2602
box -100 -472 100 472
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_0
timestamp 1666464484
transform 1 0 606 0 1 6115
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_1
timestamp 1666464484
transform 1 0 1123 0 1 4515
box 0 0 1 1
use M3_M24310590878171_256x8m81  M3_M24310590878171_256x8m81_2
timestamp 1666464484
transform 1 0 106 0 1 4515
box 0 0 1 1
use M3_M24310590878196_256x8m81  M3_M24310590878196_256x8m81_0
timestamp 1666464484
transform 1 0 606 0 1 3609
box -100 -410 100 410
<< properties >>
string GDS_END 1886982
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1886504
string path 5.615 28.025 5.615 10.575 
<< end >>
