magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 1318 89 1389
rect -31 -71 89 -1
use nmos_5p043105899832100_64x8m81  nmos_5p043105899832100_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 208 1362
<< properties >>
string GDS_END 1258766
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1258516
<< end >>
