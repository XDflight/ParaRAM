magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 5686 870
rect -86 352 1291 377
rect 1974 352 2726 377
rect 3918 352 5686 377
<< pwell >>
rect 1291 352 1974 377
rect 2726 352 3918 377
rect -86 -86 5686 352
<< mvnmos >>
rect 124 156 244 228
rect 348 156 468 228
rect 516 156 636 228
rect 740 156 860 228
rect 908 156 1028 228
rect 1185 135 1305 228
rect 1648 139 1768 232
rect 2060 124 2180 196
rect 2284 124 2404 196
rect 2452 124 2572 196
rect 2620 124 2740 196
rect 2959 185 3079 257
rect 3127 185 3247 257
rect 3351 185 3471 257
rect 3576 185 3696 257
rect 4066 156 4186 228
rect 4234 156 4354 228
rect 4458 156 4578 228
rect 4718 68 4838 232
rect 5086 68 5206 232
rect 5310 68 5430 232
<< mvpmos >>
rect 124 502 224 628
rect 348 502 448 628
rect 496 502 596 628
rect 740 502 840 628
rect 888 502 988 628
rect 1185 502 1285 687
rect 1648 497 1748 660
rect 1996 497 2096 622
rect 2236 474 2336 599
rect 2440 474 2540 599
rect 2732 497 2832 622
rect 3080 497 3180 622
rect 3372 497 3472 623
rect 3576 497 3676 623
rect 3780 497 3880 623
rect 4168 527 4268 653
rect 4372 527 4472 653
rect 4612 472 4712 716
rect 4824 472 4924 716
rect 5078 472 5178 716
rect 5282 472 5382 716
<< mvndiff >>
rect 1365 244 1437 257
rect 1365 228 1378 244
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 228
rect 636 215 740 228
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 228
rect 1028 194 1185 228
rect 1028 156 1110 194
rect 1097 148 1110 156
rect 1156 148 1185 194
rect 1097 135 1185 148
rect 1305 198 1378 228
rect 1424 198 1437 244
rect 1828 244 1900 257
rect 1828 232 1841 244
rect 1305 135 1437 198
rect 1560 198 1648 232
rect 1560 152 1573 198
rect 1619 152 1648 198
rect 1560 139 1648 152
rect 1768 198 1841 232
rect 1887 198 1900 244
rect 1768 139 1900 198
rect 2800 196 2959 257
rect 1972 183 2060 196
rect 1972 137 1985 183
rect 2031 137 2060 183
rect 1972 124 2060 137
rect 2180 183 2284 196
rect 2180 137 2209 183
rect 2255 137 2284 183
rect 2180 124 2284 137
rect 2404 124 2452 196
rect 2572 124 2620 196
rect 2740 185 2959 196
rect 3079 185 3127 257
rect 3247 244 3351 257
rect 3247 198 3276 244
rect 3322 198 3351 244
rect 3247 185 3351 198
rect 3471 244 3576 257
rect 3471 198 3500 244
rect 3546 198 3576 244
rect 3471 185 3576 198
rect 3696 244 3784 257
rect 3696 198 3725 244
rect 3771 198 3784 244
rect 4638 228 4718 232
rect 3696 185 3784 198
rect 3978 215 4066 228
rect 2740 183 2899 185
rect 2740 137 2769 183
rect 2815 137 2899 183
rect 3978 169 3991 215
rect 4037 169 4066 215
rect 3978 156 4066 169
rect 4186 156 4234 228
rect 4354 215 4458 228
rect 4354 169 4383 215
rect 4429 169 4458 215
rect 4354 156 4458 169
rect 4578 156 4718 228
rect 2740 124 2899 137
rect 4638 68 4718 156
rect 4838 187 4926 232
rect 4838 141 4867 187
rect 4913 141 4926 187
rect 4838 68 4926 141
rect 4998 143 5086 232
rect 4998 97 5011 143
rect 5057 97 5086 143
rect 4998 68 5086 97
rect 5206 209 5310 232
rect 5206 163 5235 209
rect 5281 163 5310 209
rect 5206 68 5310 163
rect 5430 143 5518 232
rect 5430 97 5459 143
rect 5505 97 5518 143
rect 5430 68 5518 97
<< mvpdiff >>
rect 1516 716 1588 729
rect 1048 634 1185 687
rect 1048 628 1075 634
rect 36 585 124 628
rect 36 539 49 585
rect 95 539 124 585
rect 36 502 124 539
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 502 348 569
rect 448 502 496 628
rect 596 595 740 628
rect 596 549 665 595
rect 711 549 740 595
rect 596 502 740 549
rect 840 502 888 628
rect 988 588 1075 628
rect 1121 588 1185 634
rect 988 502 1185 588
rect 1285 561 1393 687
rect 1285 515 1322 561
rect 1368 515 1393 561
rect 1285 502 1393 515
rect 1516 670 1529 716
rect 1575 670 1588 716
rect 1516 660 1588 670
rect 1516 497 1648 660
rect 1748 559 1836 660
rect 2600 735 2672 748
rect 2600 689 2613 735
rect 2659 689 2672 735
rect 1748 513 1777 559
rect 1823 513 1836 559
rect 1748 497 1836 513
rect 1908 571 1996 622
rect 1908 525 1921 571
rect 1967 525 1996 571
rect 1908 497 1996 525
rect 2096 599 2176 622
rect 2600 622 2672 689
rect 3240 735 3312 748
rect 3240 689 3253 735
rect 3299 689 3312 735
rect 3240 623 3312 689
rect 4532 653 4612 716
rect 4080 640 4168 653
rect 3240 622 3372 623
rect 2600 599 2732 622
rect 2096 562 2236 599
rect 2096 516 2160 562
rect 2206 516 2236 562
rect 2096 497 2236 516
rect 2156 474 2236 497
rect 2336 555 2440 599
rect 2336 509 2365 555
rect 2411 509 2440 555
rect 2336 474 2440 509
rect 2540 497 2732 599
rect 2832 556 2920 622
rect 2832 510 2861 556
rect 2907 510 2920 556
rect 2832 497 2920 510
rect 2992 556 3080 622
rect 2992 510 3005 556
rect 3051 510 3080 556
rect 2992 497 3080 510
rect 3180 497 3372 622
rect 3472 556 3576 623
rect 3472 510 3501 556
rect 3547 510 3576 556
rect 3472 497 3576 510
rect 3676 575 3780 623
rect 3676 529 3705 575
rect 3751 529 3780 575
rect 3676 497 3780 529
rect 3880 556 3976 623
rect 3880 510 3909 556
rect 3955 510 3976 556
rect 4080 594 4093 640
rect 4139 594 4168 640
rect 4080 527 4168 594
rect 4268 586 4372 653
rect 4268 540 4297 586
rect 4343 540 4372 586
rect 4268 527 4372 540
rect 4472 640 4612 653
rect 4472 594 4537 640
rect 4583 594 4612 640
rect 4472 527 4612 594
rect 3880 497 3976 510
rect 2540 474 2630 497
rect 4532 472 4612 527
rect 4712 586 4824 716
rect 4712 540 4749 586
rect 4795 540 4824 586
rect 4712 472 4824 540
rect 4924 665 5078 716
rect 4924 525 4977 665
rect 5023 525 5078 665
rect 4924 472 5078 525
rect 5178 665 5282 716
rect 5178 525 5207 665
rect 5253 525 5282 665
rect 5178 472 5282 525
rect 5382 665 5470 716
rect 5382 619 5411 665
rect 5457 619 5470 665
rect 5382 472 5470 619
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1110 148 1156 194
rect 1378 198 1424 244
rect 1573 152 1619 198
rect 1841 198 1887 244
rect 1985 137 2031 183
rect 2209 137 2255 183
rect 3276 198 3322 244
rect 3500 198 3546 244
rect 3725 198 3771 244
rect 2769 137 2815 183
rect 3991 169 4037 215
rect 4383 169 4429 215
rect 4867 141 4913 187
rect 5011 97 5057 143
rect 5235 163 5281 209
rect 5459 97 5505 143
<< mvpdiffc >>
rect 49 539 95 585
rect 263 569 309 615
rect 665 549 711 595
rect 1075 588 1121 634
rect 1322 515 1368 561
rect 1529 670 1575 716
rect 2613 689 2659 735
rect 1777 513 1823 559
rect 1921 525 1967 571
rect 3253 689 3299 735
rect 2160 516 2206 562
rect 2365 509 2411 555
rect 2861 510 2907 556
rect 3005 510 3051 556
rect 3501 510 3547 556
rect 3705 529 3751 575
rect 3909 510 3955 556
rect 4093 594 4139 640
rect 4297 540 4343 586
rect 4537 594 4583 640
rect 4749 540 4795 586
rect 4977 525 5023 665
rect 5207 525 5253 665
rect 5411 619 5457 665
<< polysilicon >>
rect 124 720 988 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 740 628 840 672
rect 888 628 988 720
rect 1185 687 1285 731
rect 1648 720 2336 760
rect 1648 660 1748 720
rect 2236 678 2336 720
rect 124 432 224 502
rect 124 351 244 432
rect 124 305 151 351
rect 197 305 244 351
rect 124 228 244 305
rect 348 351 448 502
rect 496 469 596 502
rect 496 423 525 469
rect 571 423 596 469
rect 496 410 596 423
rect 348 305 375 351
rect 421 305 448 351
rect 348 272 448 305
rect 740 407 840 502
rect 888 458 988 502
rect 740 361 753 407
rect 799 361 840 407
rect 1185 415 1285 502
rect 1996 622 2096 666
rect 2236 632 2264 678
rect 2310 632 2336 678
rect 2236 599 2336 632
rect 2440 599 2540 644
rect 2732 622 2832 666
rect 3080 622 3180 666
rect 3372 720 4268 760
rect 3372 623 3472 720
rect 3576 623 3676 667
rect 3780 623 3880 667
rect 4168 653 4268 720
rect 4612 716 4712 760
rect 4824 716 4924 760
rect 5078 716 5178 760
rect 5282 716 5382 760
rect 4372 653 4472 704
rect 1185 369 1213 415
rect 1259 413 1285 415
rect 1648 448 1748 497
rect 1259 369 1305 413
rect 740 272 840 361
rect 908 335 1028 363
rect 908 289 926 335
rect 972 289 1028 335
rect 348 228 468 272
rect 516 228 636 272
rect 740 228 860 272
rect 908 228 1028 289
rect 1185 228 1305 369
rect 1648 402 1661 448
rect 1707 402 1748 448
rect 1648 277 1748 402
rect 1996 407 2096 497
rect 2236 430 2336 474
rect 2440 430 2540 474
rect 1996 361 2009 407
rect 2055 376 2096 407
rect 2452 384 2540 430
rect 2055 361 2404 376
rect 1996 336 2404 361
rect 2284 324 2404 336
rect 2284 278 2325 324
rect 2371 278 2404 324
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1648 232 1768 277
rect 2060 196 2180 240
rect 2284 196 2404 278
rect 2452 367 2572 384
rect 2452 321 2490 367
rect 2536 321 2572 367
rect 2732 357 2832 497
rect 3080 459 3180 497
rect 3080 437 3106 459
rect 2452 196 2572 321
rect 2620 317 2832 357
rect 3007 413 3106 437
rect 3152 413 3180 459
rect 3372 437 3472 497
rect 3007 397 3180 413
rect 3228 397 3472 437
rect 3576 464 3676 497
rect 3576 418 3609 464
rect 3655 418 3676 464
rect 3780 431 3880 497
rect 4168 483 4268 527
rect 4168 466 4246 483
rect 2620 196 2740 317
rect 3007 301 3079 397
rect 3228 353 3300 397
rect 3200 317 3300 353
rect 3351 336 3471 349
rect 3200 301 3247 317
rect 2959 257 3079 301
rect 3127 257 3247 301
rect 3351 290 3388 336
rect 3434 290 3471 336
rect 3351 257 3471 290
rect 3576 301 3676 418
rect 3840 361 3880 431
rect 4108 426 4246 466
rect 4108 383 4186 426
rect 3840 340 3948 361
rect 3576 257 3696 301
rect 3840 294 3889 340
rect 3935 294 3948 340
rect 3840 281 3948 294
rect 4108 337 4121 383
rect 4167 337 4186 383
rect 4372 419 4472 527
rect 4372 378 4402 419
rect 4108 272 4186 337
rect 1185 91 1305 135
rect 124 24 636 64
rect 1648 64 1768 139
rect 4066 228 4186 272
rect 4234 373 4402 378
rect 4448 373 4472 419
rect 4612 414 4712 472
rect 4612 412 4625 414
rect 4234 338 4472 373
rect 4538 368 4625 412
rect 4671 368 4712 414
rect 4824 439 4924 472
rect 4824 412 4852 439
rect 4538 355 4712 368
rect 4798 393 4852 412
rect 4898 393 4924 439
rect 5078 416 5178 472
rect 4798 372 4924 393
rect 5086 414 5178 416
rect 4234 228 4354 338
rect 4538 272 4578 355
rect 4798 293 4838 372
rect 4458 228 4578 272
rect 4718 232 4838 293
rect 5086 368 5109 414
rect 5155 394 5178 414
rect 5282 414 5382 472
rect 5282 394 5300 414
rect 5155 368 5300 394
rect 5346 368 5382 414
rect 5086 348 5382 368
rect 5086 232 5206 348
rect 5310 288 5382 348
rect 5310 232 5430 288
rect 2959 141 3079 185
rect 3127 141 3247 185
rect 3351 141 3471 185
rect 3576 141 3696 185
rect 2060 64 2180 124
rect 2284 80 2404 124
rect 2452 80 2572 124
rect 1648 24 2180 64
rect 2620 64 2740 124
rect 4066 112 4186 156
rect 4234 112 4354 156
rect 4458 64 4578 156
rect 2620 24 4578 64
rect 4718 24 4838 68
rect 5086 24 5206 68
rect 5310 24 5430 68
<< polycontact >>
rect 151 305 197 351
rect 525 423 571 469
rect 375 305 421 351
rect 753 361 799 407
rect 2264 632 2310 678
rect 1213 369 1259 415
rect 926 289 972 335
rect 1661 402 1707 448
rect 2009 361 2055 407
rect 2325 278 2371 324
rect 2490 321 2536 367
rect 3106 413 3152 459
rect 3609 418 3655 464
rect 3388 290 3434 336
rect 3889 294 3935 340
rect 4121 337 4167 383
rect 4402 373 4448 419
rect 4625 368 4671 414
rect 4852 393 4898 439
rect 5109 368 5155 414
rect 5300 368 5346 414
<< metal1 >>
rect 0 735 5600 844
rect 0 724 2613 735
rect 252 615 320 724
rect 49 585 95 608
rect 252 569 263 615
rect 309 569 320 615
rect 1075 634 1121 724
rect 1518 716 1586 724
rect 654 549 665 595
rect 711 549 824 595
rect 1075 577 1121 588
rect 1217 632 1472 678
rect 1518 670 1529 716
rect 1575 670 1586 716
rect 2602 689 2613 724
rect 2659 724 3253 735
rect 2659 689 2670 724
rect 3240 689 3253 724
rect 3299 724 5600 735
rect 3299 689 3312 724
rect 49 523 95 539
rect 778 531 824 549
rect 1217 531 1263 632
rect 1426 624 1472 632
rect 1641 632 1967 678
rect 2253 632 2264 678
rect 2310 643 2556 678
rect 2716 643 3194 678
rect 3358 643 3655 678
rect 2310 632 3655 643
rect 1641 624 1687 632
rect 1426 578 1687 624
rect 49 477 571 523
rect 778 484 1263 531
rect 1322 561 1368 578
rect 1777 559 1823 578
rect 1368 515 1707 524
rect 1322 477 1707 515
rect 49 215 95 477
rect 525 469 571 477
rect 49 156 95 169
rect 141 351 206 430
rect 141 305 151 351
rect 197 305 206 351
rect 141 119 206 305
rect 365 351 430 430
rect 365 305 375 351
rect 421 305 430 351
rect 273 215 319 228
rect 273 60 319 169
rect 365 119 430 305
rect 525 307 571 423
rect 682 407 878 431
rect 682 361 753 407
rect 799 361 878 407
rect 682 353 878 361
rect 1026 415 1326 431
rect 1026 369 1213 415
rect 1259 369 1326 415
rect 1026 353 1326 369
rect 926 335 972 350
rect 525 289 926 307
rect 525 261 972 289
rect 1018 252 1248 298
rect 1389 255 1435 477
rect 1661 448 1707 477
rect 1661 382 1707 402
rect 1777 407 1823 513
rect 1921 571 1967 632
rect 2510 597 2762 632
rect 3148 597 3404 632
rect 1921 497 1967 525
rect 2160 562 2206 574
rect 2160 459 2206 516
rect 2336 509 2365 555
rect 2411 551 2440 555
rect 2832 551 2861 556
rect 2411 510 2861 551
rect 2907 510 2920 556
rect 2411 509 2920 510
rect 2336 505 2920 509
rect 2992 510 3005 556
rect 3051 551 3080 556
rect 3472 551 3501 556
rect 3051 510 3501 551
rect 3547 510 3558 556
rect 2992 505 3558 510
rect 2160 413 3106 459
rect 3152 413 3181 459
rect 1777 361 2009 407
rect 2055 361 2078 407
rect 1777 360 2078 361
rect 1018 215 1064 252
rect 650 169 665 215
rect 711 169 1064 215
rect 1110 194 1156 205
rect 1110 60 1156 148
rect 1202 152 1248 252
rect 1367 244 1435 255
rect 1367 198 1378 244
rect 1424 198 1435 244
rect 1481 259 1736 306
rect 1481 152 1527 259
rect 1202 106 1527 152
rect 1573 198 1619 209
rect 1573 60 1619 152
rect 1690 152 1736 259
rect 1830 244 1898 360
rect 1830 198 1841 244
rect 1887 198 1898 244
rect 1985 183 2031 196
rect 1690 137 1985 152
rect 1690 106 2031 137
rect 2209 183 2255 413
rect 3265 367 3333 505
rect 3609 464 3655 632
rect 3609 407 3655 418
rect 3705 632 4047 678
rect 3705 575 3751 632
rect 2325 324 2371 340
rect 2459 321 2490 367
rect 2536 321 3333 367
rect 3705 361 3751 529
rect 3909 556 3955 567
rect 3909 445 3955 510
rect 4001 537 4047 632
rect 4093 640 4139 724
rect 4093 583 4139 594
rect 4185 632 4463 678
rect 4185 537 4231 632
rect 4001 491 4231 537
rect 4286 540 4297 586
rect 4343 540 4354 586
rect 2325 275 2371 278
rect 2325 229 2920 275
rect 2209 124 2255 137
rect 2756 137 2769 183
rect 2815 137 2828 183
rect 2756 60 2828 137
rect 2874 152 2920 229
rect 3265 244 3333 321
rect 3265 198 3276 244
rect 3322 198 3333 244
rect 3388 336 3434 349
rect 3388 152 3434 290
rect 3489 315 3751 361
rect 3797 399 4037 445
rect 3489 244 3557 315
rect 3797 244 3843 399
rect 3489 198 3500 244
rect 3546 198 3557 244
rect 3714 198 3725 244
rect 3771 198 3843 244
rect 3889 340 3935 353
rect 3889 152 3935 294
rect 2874 106 3935 152
rect 3991 215 4037 399
rect 4121 383 4228 438
rect 4286 431 4354 540
rect 4416 548 4463 632
rect 4526 640 4594 724
rect 4526 594 4537 640
rect 4583 594 4594 640
rect 4640 632 4898 678
rect 4640 548 4686 632
rect 4416 502 4686 548
rect 4738 540 4749 586
rect 4795 540 4806 586
rect 4167 337 4228 383
rect 4121 242 4228 337
rect 4280 385 4354 431
rect 4402 419 4448 440
rect 4280 192 4326 385
rect 4402 307 4448 373
rect 4498 414 4686 431
rect 4498 368 4625 414
rect 4671 368 4686 414
rect 4498 353 4686 368
rect 4738 307 4806 540
rect 4852 439 4898 632
rect 4977 665 5023 724
rect 4977 506 5023 525
rect 5170 665 5260 676
rect 5170 525 5207 665
rect 5253 532 5260 665
rect 5411 665 5457 724
rect 5411 588 5457 619
rect 5253 525 5462 532
rect 5170 477 5462 525
rect 4852 382 4898 393
rect 4989 414 5358 419
rect 4989 368 5109 414
rect 5155 368 5300 414
rect 5346 368 5358 414
rect 4989 365 5358 368
rect 4989 307 5035 365
rect 5405 307 5462 477
rect 4402 261 5035 307
rect 4037 169 4326 192
rect 3991 143 4326 169
rect 4372 169 4383 215
rect 4429 169 4440 215
rect 4372 60 4440 169
rect 4867 187 4913 261
rect 5170 242 5462 307
rect 5170 209 5287 242
rect 4867 128 4913 141
rect 5011 143 5057 170
rect 5170 163 5235 209
rect 5281 163 5287 209
rect 5170 122 5287 163
rect 5459 143 5505 170
rect 5011 60 5057 97
rect 5459 60 5505 97
rect 0 -60 5600 60
<< labels >>
flabel metal1 s 5170 532 5260 676 0 FreeSans 400 0 0 0 Q
port 7 nsew default output
flabel metal1 s 4498 353 4686 431 0 FreeSans 400 0 0 0 RN
port 2 nsew default input
flabel metal1 s 141 119 206 430 0 FreeSans 400 0 0 0 SE
port 3 nsew default input
flabel metal1 s 4121 242 4228 438 0 FreeSans 400 0 0 0 SETN
port 4 nsew default input
flabel metal1 s 365 119 430 430 0 FreeSans 400 0 0 0 SI
port 5 nsew default input
flabel metal1 s 0 724 5600 844 0 FreeSans 400 0 0 0 VDD
port 8 nsew power bidirectional abutment
flabel metal1 s 273 215 319 228 0 FreeSans 400 0 0 0 VSS
port 11 nsew ground bidirectional abutment
flabel metal1 s 1026 353 1326 431 0 FreeSans 400 0 0 0 CLK
port 6 nsew clock input
flabel metal1 s 682 353 878 431 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 5170 477 5462 532 1 Q
port 7 nsew default output
rlabel metal1 s 5405 307 5462 477 1 Q
port 7 nsew default output
rlabel metal1 s 5170 242 5462 307 1 Q
port 7 nsew default output
rlabel metal1 s 5170 122 5287 242 1 Q
port 7 nsew default output
rlabel metal1 s 5411 689 5457 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 689 5023 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 689 4594 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 689 4139 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 3240 689 3312 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 2602 689 2670 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1518 689 1586 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 689 1121 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 689 320 724 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5411 670 5457 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 670 5023 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 670 4594 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 670 4139 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1518 670 1586 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 670 1121 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 689 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5411 594 5457 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 594 5023 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4526 594 4594 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 594 4139 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 594 1121 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 594 320 670 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 5411 588 5457 594 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 588 5023 594 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 588 4139 594 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 588 1121 594 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 588 320 594 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 583 5023 588 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4093 583 4139 588 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 583 1121 588 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 583 320 588 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 577 5023 583 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 1075 577 1121 583 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 577 320 583 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 569 5023 577 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 577 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4977 506 5023 569 1 VDD
port 8 nsew power bidirectional abutment
rlabel metal1 s 4372 209 4440 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 209 319 215 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 205 4440 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 205 1619 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 205 319 209 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 183 4440 205 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 183 1619 205 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 183 1156 205 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 205 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 170 4440 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2756 170 2828 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 170 1619 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 170 1156 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 170 319 183 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5459 60 5505 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 5011 60 5057 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 4372 60 4440 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 2756 60 2828 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1573 60 1619 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 1110 60 1156 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 170 1 VSS
port 9 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5600 60 1 VSS
port 9 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5600 784
string GDS_END 263030
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 250952
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
