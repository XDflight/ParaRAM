magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -144 -2599 1106 -2144
<< nmos >>
rect 198 -6607 318 -5245
rect 422 -6607 542 -5245
rect 644 -6607 764 -5245
<< ndiff >>
rect 78 -5291 198 -5245
rect 78 -5337 122 -5291
rect 168 -5337 198 -5291
rect 78 -5459 198 -5337
rect 78 -5505 122 -5459
rect 168 -5505 198 -5459
rect 78 -5627 198 -5505
rect 78 -5673 122 -5627
rect 168 -5673 198 -5627
rect 78 -5794 198 -5673
rect 78 -5840 122 -5794
rect 168 -5840 198 -5794
rect 78 -5962 198 -5840
rect 78 -6008 122 -5962
rect 168 -6008 198 -5962
rect 78 -6130 198 -6008
rect 78 -6176 122 -6130
rect 168 -6176 198 -6130
rect 78 -6298 198 -6176
rect 78 -6344 122 -6298
rect 168 -6344 198 -6298
rect 78 -6465 198 -6344
rect 78 -6511 122 -6465
rect 168 -6511 198 -6465
rect 78 -6607 198 -6511
rect 318 -6607 422 -5245
rect 542 -6607 644 -5245
rect 764 -5291 883 -5245
rect 764 -5337 794 -5291
rect 840 -5337 883 -5291
rect 764 -5459 883 -5337
rect 764 -5505 794 -5459
rect 840 -5505 883 -5459
rect 764 -5627 883 -5505
rect 764 -5673 794 -5627
rect 840 -5673 883 -5627
rect 764 -5794 883 -5673
rect 764 -5840 794 -5794
rect 840 -5840 883 -5794
rect 764 -5962 883 -5840
rect 764 -6008 794 -5962
rect 840 -6008 883 -5962
rect 764 -6130 883 -6008
rect 764 -6176 794 -6130
rect 840 -6176 883 -6130
rect 764 -6298 883 -6176
rect 764 -6344 794 -6298
rect 840 -6344 883 -6298
rect 764 -6465 883 -6344
rect 764 -6511 794 -6465
rect 840 -6511 883 -6465
rect 764 -6607 883 -6511
<< ndiffc >>
rect 122 -5337 168 -5291
rect 122 -5505 168 -5459
rect 122 -5673 168 -5627
rect 122 -5840 168 -5794
rect 122 -6008 168 -5962
rect 122 -6176 168 -6130
rect 122 -6344 168 -6298
rect 122 -6511 168 -6465
rect 794 -5337 840 -5291
rect 794 -5505 840 -5459
rect 794 -5673 840 -5627
rect 794 -5840 840 -5794
rect 794 -6008 840 -5962
rect 794 -6176 840 -6130
rect 794 -6344 840 -6298
rect 794 -6511 840 -6465
<< psubdiff >>
rect -1 186 963 245
rect -1 140 212 186
rect 258 140 370 186
rect 416 140 528 186
rect 574 140 686 186
rect 732 140 963 186
rect -1 81 963 140
rect -1 -6883 963 -6823
rect -1 -6929 212 -6883
rect 258 -6929 370 -6883
rect 416 -6929 528 -6883
rect 574 -6929 686 -6883
rect 732 -6929 963 -6883
rect -1 -6988 963 -6929
<< nsubdiff >>
rect -1 -2349 963 -2292
rect -1 -2395 201 -2349
rect 247 -2395 359 -2349
rect 405 -2395 517 -2349
rect 563 -2395 963 -2349
rect -1 -2452 963 -2395
<< psubdiffcont >>
rect 212 140 258 186
rect 370 140 416 186
rect 528 140 574 186
rect 686 140 732 186
rect 212 -6929 258 -6883
rect 370 -6929 416 -6883
rect 528 -6929 574 -6883
rect 686 -6929 732 -6883
<< nsubdiffcont >>
rect 201 -2395 247 -2349
rect 359 -2395 405 -2349
rect 517 -2395 563 -2349
<< polysilicon >>
rect 197 -662 317 -620
rect 421 -662 541 -620
rect 645 -662 765 -620
rect 197 -799 765 -662
rect 197 -858 317 -799
rect 421 -858 541 -799
rect 645 -858 765 -799
rect 197 -2094 317 -2048
rect 421 -2094 541 -2038
rect 645 -2094 765 -2048
rect 197 -2113 765 -2094
rect 197 -2159 378 -2113
rect 612 -2159 765 -2113
rect 197 -2178 765 -2159
rect 198 -4377 316 -3911
rect 421 -4224 541 -3911
rect 645 -4077 765 -3911
rect 421 -4311 542 -4224
rect 198 -4515 317 -4377
rect 198 -4982 318 -4515
rect 197 -5120 318 -4982
rect 198 -5245 318 -5120
rect 422 -5245 542 -4311
rect 645 -4579 764 -4077
rect 644 -5245 764 -4579
rect 198 -6680 318 -6607
rect 422 -6680 542 -6607
rect 644 -6680 764 -6607
<< polycontact >>
rect 378 -2159 612 -2113
<< metal1 >>
rect -1 186 963 237
rect -1 167 212 186
rect -1 115 119 167
rect 171 140 212 167
rect 258 140 370 186
rect 416 140 528 186
rect 574 167 686 186
rect 619 140 686 167
rect 732 140 963 186
rect 171 115 567 140
rect 619 115 963 140
rect -1 -51 963 115
rect -1 -55 119 -51
rect 81 -103 119 -55
rect 171 -55 567 -51
rect 171 -103 209 -55
rect 81 -269 209 -103
rect 529 -103 567 -55
rect 619 -55 963 -51
rect 619 -103 657 -55
rect 81 -321 119 -269
rect 171 -321 209 -269
rect 81 -487 209 -321
rect 81 -539 119 -487
rect 171 -539 209 -487
rect 81 -579 209 -539
rect 303 -184 431 -145
rect 303 -236 341 -184
rect 393 -236 431 -184
rect 303 -402 431 -236
rect 303 -454 341 -402
rect 393 -454 431 -402
rect 303 -620 431 -454
rect 529 -269 657 -103
rect 529 -321 567 -269
rect 619 -321 657 -269
rect 529 -487 657 -321
rect 529 -539 567 -487
rect 619 -539 657 -487
rect 529 -579 657 -539
rect 303 -672 341 -620
rect 393 -666 431 -620
rect 759 -666 874 -507
rect 393 -672 874 -666
rect 303 -712 874 -672
rect 311 -713 874 -712
rect 312 -785 874 -713
rect 312 -786 427 -785
rect 312 -930 426 -786
rect 759 -930 874 -785
rect 81 -1338 209 -1299
rect 81 -1390 119 -1338
rect 171 -1390 209 -1338
rect 81 -1556 209 -1390
rect 81 -1608 119 -1556
rect 171 -1608 209 -1556
rect 81 -1774 209 -1608
rect 81 -1826 119 -1774
rect 171 -1826 209 -1774
rect 81 -1866 209 -1826
rect 529 -1338 657 -1299
rect 529 -1390 567 -1338
rect 619 -1390 657 -1338
rect 529 -1556 657 -1390
rect 529 -1608 567 -1556
rect 619 -1608 657 -1556
rect 529 -1774 657 -1608
rect 529 -1826 567 -1774
rect 619 -1826 657 -1774
rect 529 -1866 657 -1826
rect 200 -2113 874 -2076
rect 200 -2159 378 -2113
rect 612 -2159 874 -2113
rect 200 -2195 874 -2159
rect -1 -2349 650 -2312
rect -1 -2395 201 -2349
rect 247 -2395 359 -2349
rect 405 -2395 517 -2349
rect 563 -2395 650 -2349
rect -1 -2407 650 -2395
rect -1 -2431 652 -2407
rect 81 -2447 209 -2431
rect 81 -2499 119 -2447
rect 171 -2499 209 -2447
rect 81 -2665 209 -2499
rect 81 -2717 119 -2665
rect 171 -2717 209 -2665
rect 81 -2882 209 -2717
rect 81 -2934 119 -2882
rect 171 -2934 209 -2882
rect 81 -3100 209 -2934
rect 81 -3152 119 -3100
rect 171 -3152 209 -3100
rect 81 -3318 209 -3152
rect 81 -3370 119 -3318
rect 171 -3370 209 -3318
rect 81 -3535 209 -3370
rect 525 -2448 652 -2431
rect 525 -2500 563 -2448
rect 615 -2500 652 -2448
rect 525 -2665 652 -2500
rect 525 -2717 563 -2665
rect 615 -2717 652 -2665
rect 525 -2883 652 -2717
rect 759 -2771 874 -2195
rect 525 -2935 563 -2883
rect 615 -2935 652 -2883
rect 525 -3101 652 -2935
rect 525 -3153 563 -3101
rect 615 -3153 652 -3101
rect 525 -3318 652 -3153
rect 525 -3370 563 -3318
rect 615 -3370 652 -3318
rect 525 -3411 652 -3370
rect 81 -3587 119 -3535
rect 171 -3587 209 -3535
rect 81 -3753 209 -3587
rect 81 -3805 119 -3753
rect 171 -3805 209 -3753
rect 81 -3845 209 -3805
rect 94 -3846 209 -3845
rect 307 -3553 431 -3513
rect 307 -3605 343 -3553
rect 395 -3605 431 -3553
rect 307 -3771 431 -3605
rect 307 -3823 343 -3771
rect 395 -3823 431 -3771
rect 307 -3863 431 -3823
rect 755 -3553 879 -3513
rect 755 -3605 791 -3553
rect 843 -3605 879 -3553
rect 755 -3771 879 -3605
rect 755 -3823 791 -3771
rect 843 -3823 879 -3771
rect 755 -3863 879 -3823
rect -58 -4088 1020 -3996
rect -58 -4290 1020 -4198
rect -58 -4492 1020 -4400
rect -58 -4694 1020 -4602
rect -58 -4895 1020 -4803
rect -58 -5097 1020 -5005
rect 88 -5291 202 -5254
rect 88 -5337 122 -5291
rect 168 -5337 202 -5291
rect 88 -5350 202 -5337
rect 759 -5291 874 -5254
rect 759 -5337 794 -5291
rect 840 -5337 874 -5291
rect 87 -5459 203 -5350
rect 759 -5404 874 -5337
rect 87 -5505 122 -5459
rect 168 -5505 203 -5459
rect 87 -5627 203 -5505
rect 87 -5673 122 -5627
rect 168 -5673 203 -5627
rect 87 -5794 203 -5673
rect 87 -5840 122 -5794
rect 168 -5840 203 -5794
rect 87 -5962 203 -5840
rect 87 -6008 122 -5962
rect 168 -6008 203 -5962
rect 87 -6130 203 -6008
rect 87 -6176 122 -6130
rect 168 -6176 203 -6130
rect 87 -6298 203 -6176
rect 87 -6344 122 -6298
rect 168 -6344 203 -6298
rect 87 -6465 203 -6344
rect 753 -5445 880 -5404
rect 753 -5497 791 -5445
rect 843 -5497 880 -5445
rect 753 -5505 794 -5497
rect 840 -5505 880 -5497
rect 753 -5627 880 -5505
rect 753 -5662 794 -5627
rect 840 -5662 880 -5627
rect 753 -5714 791 -5662
rect 843 -5714 880 -5662
rect 753 -5794 880 -5714
rect 753 -5840 794 -5794
rect 840 -5840 880 -5794
rect 753 -5880 880 -5840
rect 753 -5932 791 -5880
rect 843 -5932 880 -5880
rect 753 -5962 880 -5932
rect 753 -6008 794 -5962
rect 840 -6008 880 -5962
rect 753 -6098 880 -6008
rect 753 -6150 791 -6098
rect 843 -6150 880 -6098
rect 753 -6176 794 -6150
rect 840 -6176 880 -6150
rect 753 -6298 880 -6176
rect 753 -6315 794 -6298
rect 840 -6315 880 -6298
rect 753 -6367 791 -6315
rect 843 -6367 880 -6315
rect 753 -6408 880 -6367
rect 87 -6511 122 -6465
rect 168 -6511 203 -6465
rect 87 -6687 203 -6511
rect 759 -6465 874 -6408
rect 759 -6511 794 -6465
rect 840 -6511 874 -6465
rect 759 -6598 874 -6511
rect 8 -6883 963 -6687
rect 8 -6929 212 -6883
rect 258 -6929 370 -6883
rect 416 -6929 528 -6883
rect 574 -6929 686 -6883
rect 732 -6929 963 -6883
rect 8 -6979 963 -6929
<< via1 >>
rect 119 115 171 167
rect 567 140 574 167
rect 574 140 619 167
rect 567 115 619 140
rect 119 -103 171 -51
rect 567 -103 619 -51
rect 119 -321 171 -269
rect 119 -539 171 -487
rect 341 -236 393 -184
rect 341 -454 393 -402
rect 567 -321 619 -269
rect 567 -539 619 -487
rect 341 -672 393 -620
rect 119 -1390 171 -1338
rect 119 -1608 171 -1556
rect 119 -1826 171 -1774
rect 567 -1390 619 -1338
rect 567 -1608 619 -1556
rect 567 -1826 619 -1774
rect 119 -2499 171 -2447
rect 119 -2717 171 -2665
rect 119 -2934 171 -2882
rect 119 -3152 171 -3100
rect 119 -3370 171 -3318
rect 563 -2500 615 -2448
rect 563 -2717 615 -2665
rect 563 -2935 615 -2883
rect 563 -3153 615 -3101
rect 563 -3370 615 -3318
rect 119 -3587 171 -3535
rect 119 -3805 171 -3753
rect 343 -3605 395 -3553
rect 343 -3823 395 -3771
rect 791 -3605 843 -3553
rect 791 -3823 843 -3771
rect 791 -5459 843 -5445
rect 791 -5497 794 -5459
rect 794 -5497 840 -5459
rect 840 -5497 843 -5459
rect 791 -5673 794 -5662
rect 794 -5673 840 -5662
rect 840 -5673 843 -5662
rect 791 -5714 843 -5673
rect 791 -5932 843 -5880
rect 791 -6130 843 -6098
rect 791 -6150 794 -6130
rect 794 -6150 840 -6130
rect 840 -6150 843 -6130
rect 791 -6344 794 -6315
rect 794 -6344 840 -6315
rect 840 -6344 843 -6315
rect 791 -6367 843 -6344
<< metal2 >>
rect 81 169 209 206
rect 81 113 117 169
rect 173 113 209 169
rect 81 -49 209 113
rect 81 -105 117 -49
rect 173 -105 209 -49
rect 81 -267 209 -105
rect 81 -323 117 -267
rect 173 -323 209 -267
rect 81 -485 209 -323
rect 81 -541 117 -485
rect 173 -541 209 -485
rect 81 -579 209 -541
rect 303 -184 431 327
rect 303 -236 341 -184
rect 393 -236 431 -184
rect 303 -402 431 -236
rect 303 -454 341 -402
rect 393 -454 431 -402
rect 303 -620 431 -454
rect 529 169 657 206
rect 529 113 565 169
rect 621 113 657 169
rect 529 -49 657 113
rect 529 -105 565 -49
rect 621 -105 657 -49
rect 529 -267 657 -105
rect 529 -323 565 -267
rect 621 -323 657 -267
rect 529 -485 657 -323
rect 529 -541 565 -485
rect 621 -541 657 -485
rect 529 -579 657 -541
rect 303 -672 341 -620
rect 393 -672 431 -620
rect 303 -712 431 -672
rect 81 -1336 209 -1299
rect 81 -1392 117 -1336
rect 173 -1392 209 -1336
rect 81 -1554 209 -1392
rect 81 -1610 117 -1554
rect 173 -1610 209 -1554
rect 81 -1772 209 -1610
rect 81 -1828 117 -1772
rect 173 -1828 209 -1772
rect 81 -1866 209 -1828
rect 529 -1336 657 -1299
rect 529 -1392 565 -1336
rect 621 -1392 657 -1336
rect 529 -1554 657 -1392
rect 529 -1610 565 -1554
rect 621 -1610 657 -1554
rect 529 -1772 657 -1610
rect 529 -1828 565 -1772
rect 621 -1828 657 -1772
rect 529 -1866 657 -1828
rect 81 -2445 209 -2408
rect 81 -2501 117 -2445
rect 173 -2501 209 -2445
rect 81 -2663 209 -2501
rect 81 -2719 117 -2663
rect 173 -2719 209 -2663
rect 81 -2880 209 -2719
rect 81 -2936 117 -2880
rect 173 -2936 209 -2880
rect 81 -3098 209 -2936
rect 81 -3154 117 -3098
rect 173 -3154 209 -3098
rect 81 -3316 209 -3154
rect 81 -3372 117 -3316
rect 173 -3372 209 -3316
rect 81 -3533 209 -3372
rect 525 -2446 652 -2407
rect 525 -2502 561 -2446
rect 617 -2502 652 -2446
rect 525 -2663 652 -2502
rect 525 -2719 561 -2663
rect 617 -2719 652 -2663
rect 525 -2881 652 -2719
rect 525 -2937 561 -2881
rect 617 -2937 652 -2881
rect 525 -3099 652 -2937
rect 525 -3155 561 -3099
rect 617 -3155 652 -3099
rect 525 -3316 652 -3155
rect 525 -3372 561 -3316
rect 617 -3372 652 -3316
rect 525 -3411 652 -3372
rect 81 -3589 117 -3533
rect 173 -3589 209 -3533
rect 81 -3751 209 -3589
rect 81 -3807 117 -3751
rect 173 -3807 209 -3751
rect 81 -3845 209 -3807
rect 305 -3553 881 -3513
rect 305 -3605 343 -3553
rect 395 -3605 791 -3553
rect 843 -3605 881 -3553
rect 305 -3771 881 -3605
rect 305 -3823 343 -3771
rect 395 -3823 791 -3771
rect 843 -3823 881 -3771
rect 305 -3864 881 -3823
rect 752 -3865 881 -3864
rect 753 -5445 881 -3865
rect 753 -5497 791 -5445
rect 843 -5497 881 -5445
rect 753 -5546 881 -5497
rect 753 -5662 880 -5546
rect 753 -5714 791 -5662
rect 843 -5714 880 -5662
rect 753 -5880 880 -5714
rect 753 -5932 791 -5880
rect 843 -5932 880 -5880
rect 753 -6098 880 -5932
rect 753 -6150 791 -6098
rect 843 -6150 880 -6098
rect 753 -6315 880 -6150
rect 753 -6367 791 -6315
rect 843 -6367 880 -6315
rect 753 -6408 880 -6367
<< via2 >>
rect 117 167 173 169
rect 117 115 119 167
rect 119 115 171 167
rect 171 115 173 167
rect 117 113 173 115
rect 117 -51 173 -49
rect 117 -103 119 -51
rect 119 -103 171 -51
rect 171 -103 173 -51
rect 117 -105 173 -103
rect 117 -269 173 -267
rect 117 -321 119 -269
rect 119 -321 171 -269
rect 171 -321 173 -269
rect 117 -323 173 -321
rect 117 -487 173 -485
rect 117 -539 119 -487
rect 119 -539 171 -487
rect 171 -539 173 -487
rect 117 -541 173 -539
rect 565 167 621 169
rect 565 115 567 167
rect 567 115 619 167
rect 619 115 621 167
rect 565 113 621 115
rect 565 -51 621 -49
rect 565 -103 567 -51
rect 567 -103 619 -51
rect 619 -103 621 -51
rect 565 -105 621 -103
rect 565 -269 621 -267
rect 565 -321 567 -269
rect 567 -321 619 -269
rect 619 -321 621 -269
rect 565 -323 621 -321
rect 565 -487 621 -485
rect 565 -539 567 -487
rect 567 -539 619 -487
rect 619 -539 621 -487
rect 565 -541 621 -539
rect 117 -1338 173 -1336
rect 117 -1390 119 -1338
rect 119 -1390 171 -1338
rect 171 -1390 173 -1338
rect 117 -1392 173 -1390
rect 117 -1556 173 -1554
rect 117 -1608 119 -1556
rect 119 -1608 171 -1556
rect 171 -1608 173 -1556
rect 117 -1610 173 -1608
rect 117 -1774 173 -1772
rect 117 -1826 119 -1774
rect 119 -1826 171 -1774
rect 171 -1826 173 -1774
rect 117 -1828 173 -1826
rect 565 -1338 621 -1336
rect 565 -1390 567 -1338
rect 567 -1390 619 -1338
rect 619 -1390 621 -1338
rect 565 -1392 621 -1390
rect 565 -1556 621 -1554
rect 565 -1608 567 -1556
rect 567 -1608 619 -1556
rect 619 -1608 621 -1556
rect 565 -1610 621 -1608
rect 565 -1774 621 -1772
rect 565 -1826 567 -1774
rect 567 -1826 619 -1774
rect 619 -1826 621 -1774
rect 565 -1828 621 -1826
rect 117 -2447 173 -2445
rect 117 -2499 119 -2447
rect 119 -2499 171 -2447
rect 171 -2499 173 -2447
rect 117 -2501 173 -2499
rect 117 -2665 173 -2663
rect 117 -2717 119 -2665
rect 119 -2717 171 -2665
rect 171 -2717 173 -2665
rect 117 -2719 173 -2717
rect 117 -2882 173 -2880
rect 117 -2934 119 -2882
rect 119 -2934 171 -2882
rect 171 -2934 173 -2882
rect 117 -2936 173 -2934
rect 117 -3100 173 -3098
rect 117 -3152 119 -3100
rect 119 -3152 171 -3100
rect 171 -3152 173 -3100
rect 117 -3154 173 -3152
rect 117 -3318 173 -3316
rect 117 -3370 119 -3318
rect 119 -3370 171 -3318
rect 171 -3370 173 -3318
rect 117 -3372 173 -3370
rect 561 -2448 617 -2446
rect 561 -2500 563 -2448
rect 563 -2500 615 -2448
rect 615 -2500 617 -2448
rect 561 -2502 617 -2500
rect 561 -2665 617 -2663
rect 561 -2717 563 -2665
rect 563 -2717 615 -2665
rect 615 -2717 617 -2665
rect 561 -2719 617 -2717
rect 561 -2883 617 -2881
rect 561 -2935 563 -2883
rect 563 -2935 615 -2883
rect 615 -2935 617 -2883
rect 561 -2937 617 -2935
rect 561 -3101 617 -3099
rect 561 -3153 563 -3101
rect 563 -3153 615 -3101
rect 615 -3153 617 -3101
rect 561 -3155 617 -3153
rect 561 -3318 617 -3316
rect 561 -3370 563 -3318
rect 563 -3370 615 -3318
rect 615 -3370 617 -3318
rect 561 -3372 617 -3370
rect 117 -3535 173 -3533
rect 117 -3587 119 -3535
rect 119 -3587 171 -3535
rect 171 -3587 173 -3535
rect 117 -3589 173 -3587
rect 117 -3753 173 -3751
rect 117 -3805 119 -3753
rect 119 -3805 171 -3753
rect 171 -3805 173 -3753
rect 117 -3807 173 -3805
<< metal3 >>
rect -52 169 1106 327
rect -52 113 117 169
rect 173 113 565 169
rect 621 113 1106 169
rect -52 -49 1106 113
rect -52 -105 117 -49
rect 173 -105 565 -49
rect 621 -105 1106 -49
rect -52 -267 1106 -105
rect -52 -323 117 -267
rect 173 -323 565 -267
rect 621 -323 1106 -267
rect -52 -485 1106 -323
rect -52 -541 117 -485
rect 173 -541 565 -485
rect 621 -541 1106 -485
rect -52 -624 1106 -541
rect -58 -1336 1106 -1262
rect -58 -1392 117 -1336
rect 173 -1392 565 -1336
rect 621 -1392 1106 -1336
rect -58 -1554 1106 -1392
rect -58 -1610 117 -1554
rect 173 -1610 565 -1554
rect 621 -1610 1106 -1554
rect -58 -1772 1106 -1610
rect -58 -1828 117 -1772
rect 173 -1828 565 -1772
rect 621 -1828 1106 -1772
rect -58 -2171 1106 -1828
rect -58 -2445 919 -2171
rect -58 -2501 117 -2445
rect 173 -2446 919 -2445
rect 173 -2501 561 -2446
rect -58 -2502 561 -2501
rect 617 -2502 919 -2446
rect -58 -2663 919 -2502
rect -58 -2719 117 -2663
rect 173 -2719 561 -2663
rect 617 -2719 919 -2663
rect -58 -2880 919 -2719
rect -58 -2936 117 -2880
rect 173 -2881 919 -2880
rect 173 -2936 561 -2881
rect -58 -2937 561 -2936
rect 617 -2937 919 -2881
rect -58 -3098 919 -2937
rect -58 -3154 117 -3098
rect 173 -3099 919 -3098
rect 173 -3154 561 -3099
rect -58 -3155 561 -3154
rect 617 -3155 919 -3099
rect -58 -3316 919 -3155
rect -58 -3372 117 -3316
rect 173 -3372 561 -3316
rect 617 -3372 919 -3316
rect -58 -3533 919 -3372
rect -58 -3589 117 -3533
rect 173 -3589 919 -3533
rect -58 -3751 919 -3589
rect -58 -3807 117 -3751
rect 173 -3807 919 -3751
rect -58 -3896 919 -3807
rect -1 -7124 963 -5286
use M1_POLY24310589983234_64x8m81  M1_POLY24310589983234_64x8m81_0
timestamp 1666464484
transform 1 0 495 0 1 -2136
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1666464484
transform 1 0 369 0 1 -3688
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1666464484
transform 1 0 817 0 1 -3688
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_0
timestamp 1666464484
transform 1 0 589 0 1 -2909
box 0 0 1 1
use M2_M1$$43378732_64x8m81  M2_M1$$43378732_64x8m81_1
timestamp 1666464484
transform 1 0 817 0 1 -5906
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_0
timestamp 1666464484
transform 1 0 593 0 1 -186
box 0 0 1 1
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_1
timestamp 1666464484
transform 1 0 145 0 1 -186
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_0
timestamp 1666464484
transform 1 0 367 0 1 -428
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_1
timestamp 1666464484
transform 1 0 593 0 1 -1582
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_2
timestamp 1666464484
transform 1 0 145 0 1 -1582
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -3126
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_0
timestamp 1666464484
transform 1 0 593 0 1 -1582
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_1
timestamp 1666464484
transform 1 0 145 0 1 -1582
box 0 0 1 1
use M3_M2$$47332396_64x8m81  M3_M2$$47332396_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -3126
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -186
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_1
timestamp 1666464484
transform 1 0 593 0 1 -186
box 0 0 1 1
use M3_M2$$47819820_64x8m81  M3_M2$$47819820_64x8m81_0
timestamp 1666464484
transform 1 0 589 0 1 -2909
box 0 0 1 1
use nmos_1p2$$46551084_64x8m81  nmos_1p2$$46551084_64x8m81_0
timestamp 1666464484
transform 1 0 676 0 -1 -136
box -119 -73 177 527
use nmos_1p2$$46551084_64x8m81  nmos_1p2$$46551084_64x8m81_1
timestamp 1666464484
transform 1 0 452 0 -1 -136
box -119 -73 177 527
use nmos_1p2$$46551084_64x8m81  nmos_1p2$$46551084_64x8m81_2
timestamp 1666464484
transform 1 0 228 0 -1 -136
box -119 -73 177 527
use pmos_1p2$$47820844_64x8m81  pmos_1p2$$47820844_64x8m81_0
timestamp 1666464484
transform 1 0 228 0 -1 -871
box -286 -141 344 1275
use pmos_1p2$$47820844_64x8m81  pmos_1p2$$47820844_64x8m81_1
timestamp 1666464484
transform 1 0 676 0 -1 -871
box -286 -141 344 1275
use pmos_1p2$$47820844_64x8m81  pmos_1p2$$47820844_64x8m81_2
timestamp 1666464484
transform 1 0 452 0 -1 -871
box -286 -141 344 1275
use pmos_1p2$$47821868_64x8m81  pmos_1p2$$47821868_64x8m81_0
timestamp 1666464484
transform 1 0 228 0 1 -3872
box -286 -142 344 1275
use pmos_1p2$$47821868_64x8m81  pmos_1p2$$47821868_64x8m81_1
timestamp 1666464484
transform 1 0 452 0 1 -3872
box -286 -142 344 1275
use pmos_1p2$$47821868_64x8m81  pmos_1p2$$47821868_64x8m81_2
timestamp 1666464484
transform 1 0 676 0 1 -3872
box -286 -142 344 1275
<< properties >>
string GDS_END 392816
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 387024
<< end >>
