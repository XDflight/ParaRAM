magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 2774 870
rect -86 352 678 377
rect 1047 352 2774 377
<< pwell >>
rect 678 352 1047 377
rect -86 -86 2774 352
<< mvnmos >>
rect 124 68 244 232
rect 348 68 468 232
rect 572 68 692 232
rect 1033 68 1153 232
rect 1283 68 1403 232
rect 1507 68 1627 232
rect 1731 68 1851 232
rect 1955 68 2075 232
rect 2179 68 2299 232
rect 2403 68 2523 232
<< mvpmos >>
rect 173 497 273 716
rect 377 497 477 716
rect 581 497 681 716
rect 1053 497 1153 716
rect 1293 480 1393 716
rect 1497 480 1597 716
rect 1701 480 1801 716
rect 1905 480 2005 716
rect 2109 480 2209 716
rect 2313 480 2413 716
<< mvndiff >>
rect 752 244 824 257
rect 752 232 765 244
rect 36 192 124 232
rect 36 146 49 192
rect 95 146 124 192
rect 36 68 124 146
rect 244 139 348 232
rect 244 93 273 139
rect 319 93 348 139
rect 244 68 348 93
rect 468 166 572 232
rect 468 120 497 166
rect 543 120 572 166
rect 468 68 572 120
rect 692 198 765 232
rect 811 198 824 244
rect 692 68 824 198
rect 901 244 973 257
rect 901 198 914 244
rect 960 232 973 244
rect 960 198 1033 232
rect 901 68 1033 198
rect 1153 127 1283 232
rect 1153 81 1208 127
rect 1254 81 1283 127
rect 1153 68 1283 81
rect 1403 219 1507 232
rect 1403 173 1432 219
rect 1478 173 1507 219
rect 1403 68 1507 173
rect 1627 127 1731 232
rect 1627 81 1656 127
rect 1702 81 1731 127
rect 1627 68 1731 81
rect 1851 200 1955 232
rect 1851 154 1880 200
rect 1926 154 1955 200
rect 1851 68 1955 154
rect 2075 127 2179 232
rect 2075 81 2104 127
rect 2150 81 2179 127
rect 2075 68 2179 81
rect 2299 200 2403 232
rect 2299 154 2328 200
rect 2374 154 2403 200
rect 2299 68 2403 154
rect 2523 200 2611 232
rect 2523 154 2552 200
rect 2598 154 2611 200
rect 2523 68 2611 154
<< mvpdiff >>
rect 85 665 173 716
rect 85 525 98 665
rect 144 525 173 665
rect 85 497 173 525
rect 273 703 377 716
rect 273 657 302 703
rect 348 657 377 703
rect 273 497 377 657
rect 477 671 581 716
rect 477 625 506 671
rect 552 625 581 671
rect 477 497 581 625
rect 681 567 769 716
rect 681 521 710 567
rect 756 521 769 567
rect 681 497 769 521
rect 965 567 1053 716
rect 965 521 978 567
rect 1024 521 1053 567
rect 965 497 1053 521
rect 1153 703 1293 716
rect 1153 657 1208 703
rect 1254 657 1293 703
rect 1153 497 1293 657
rect 1213 480 1293 497
rect 1393 665 1497 716
rect 1393 525 1422 665
rect 1468 525 1497 665
rect 1393 480 1497 525
rect 1597 703 1701 716
rect 1597 563 1626 703
rect 1672 563 1701 703
rect 1597 480 1701 563
rect 1801 665 1905 716
rect 1801 525 1830 665
rect 1876 525 1905 665
rect 1801 480 1905 525
rect 2005 665 2109 716
rect 2005 619 2034 665
rect 2080 619 2109 665
rect 2005 480 2109 619
rect 2209 665 2313 716
rect 2209 525 2238 665
rect 2284 525 2313 665
rect 2209 480 2313 525
rect 2413 665 2501 716
rect 2413 525 2442 665
rect 2488 525 2501 665
rect 2413 480 2501 525
<< mvndiffc >>
rect 49 146 95 192
rect 273 93 319 139
rect 497 120 543 166
rect 765 198 811 244
rect 914 198 960 244
rect 1208 81 1254 127
rect 1432 173 1478 219
rect 1656 81 1702 127
rect 1880 154 1926 200
rect 2104 81 2150 127
rect 2328 154 2374 200
rect 2552 154 2598 200
<< mvpdiffc >>
rect 98 525 144 665
rect 302 657 348 703
rect 506 625 552 671
rect 710 521 756 567
rect 978 521 1024 567
rect 1208 657 1254 703
rect 1422 525 1468 665
rect 1626 563 1672 703
rect 1830 525 1876 665
rect 2034 619 2080 665
rect 2238 525 2284 665
rect 2442 525 2488 665
<< polysilicon >>
rect 173 716 273 760
rect 377 716 477 760
rect 581 716 681 760
rect 1053 716 1153 760
rect 1293 716 1393 760
rect 1497 716 1597 760
rect 1701 716 1801 760
rect 1905 716 2005 760
rect 2109 716 2209 760
rect 2313 716 2413 760
rect 173 412 273 497
rect 377 412 477 497
rect 581 464 681 497
rect 581 418 594 464
rect 640 418 681 464
rect 124 399 533 412
rect 581 405 681 418
rect 1053 405 1153 497
rect 124 353 172 399
rect 218 372 533 399
rect 218 353 244 372
rect 124 232 244 353
rect 493 357 533 372
rect 1053 359 1080 405
rect 1126 359 1153 405
rect 348 311 433 324
rect 493 317 612 357
rect 348 265 374 311
rect 420 276 433 311
rect 572 288 612 317
rect 420 265 468 276
rect 348 232 468 265
rect 572 232 692 288
rect 1053 287 1153 359
rect 1293 418 1393 480
rect 1497 418 1597 480
rect 1293 405 1597 418
rect 1293 359 1335 405
rect 1569 359 1597 405
rect 1701 439 1801 480
rect 1701 393 1731 439
rect 1777 420 1801 439
rect 1905 439 2005 480
rect 1905 420 1933 439
rect 1777 393 1933 420
rect 1979 420 2005 439
rect 2109 420 2209 480
rect 2313 420 2413 480
rect 1979 393 2413 420
rect 1701 380 2413 393
rect 1293 346 1597 359
rect 1293 300 1403 346
rect 1033 232 1153 287
rect 1283 232 1403 300
rect 1507 287 1597 346
rect 1731 319 2523 332
rect 1507 232 1627 287
rect 1731 273 1744 319
rect 1790 292 1968 319
rect 1790 273 1851 292
rect 1731 232 1851 273
rect 1955 273 1968 292
rect 2014 292 2523 319
rect 2014 273 2075 292
rect 1955 232 2075 273
rect 2179 232 2299 292
rect 2403 232 2523 292
rect 124 24 244 68
rect 348 24 468 68
rect 572 24 692 68
rect 1033 24 1153 68
rect 1283 24 1403 68
rect 1507 24 1627 68
rect 1731 24 1851 68
rect 1955 24 2075 68
rect 2179 24 2299 68
rect 2403 24 2523 68
<< polycontact >>
rect 594 418 640 464
rect 172 353 218 399
rect 1080 359 1126 405
rect 374 265 420 311
rect 1335 359 1569 405
rect 1731 393 1777 439
rect 1933 393 1979 439
rect 1744 273 1790 319
rect 1968 273 2014 319
<< metal1 >>
rect 0 724 2688 844
rect 291 703 359 724
rect 98 665 144 676
rect 291 657 302 703
rect 348 657 359 703
rect 1197 703 1265 724
rect 495 625 506 671
rect 552 625 1125 671
rect 1197 657 1208 703
rect 1254 657 1265 703
rect 1615 703 1683 724
rect 1422 665 1468 676
rect 802 624 1125 625
rect 709 567 756 578
rect 144 525 420 548
rect 98 502 420 525
rect 374 464 420 502
rect 709 521 710 567
rect 74 399 324 430
rect 74 353 172 399
rect 218 353 324 399
rect 74 352 324 353
rect 374 418 594 464
rect 640 418 652 464
rect 374 417 652 418
rect 374 311 420 417
rect 709 361 756 521
rect 374 245 420 265
rect 49 198 420 245
rect 595 315 756 361
rect 49 192 95 198
rect 595 177 641 315
rect 802 269 848 624
rect 1079 611 1125 624
rect 978 567 1024 578
rect 1079 565 1422 611
rect 978 519 1024 521
rect 1615 563 1626 703
rect 1672 563 1683 703
rect 1822 665 1882 676
rect 978 473 1366 519
rect 895 405 1214 427
rect 895 359 1080 405
rect 1126 359 1214 405
rect 895 358 1214 359
rect 1320 425 1366 473
rect 1422 517 1468 525
rect 1822 525 1830 665
rect 1876 532 1882 665
rect 2034 665 2080 724
rect 2034 604 2080 619
rect 2238 665 2284 676
rect 1876 525 2238 532
rect 1422 471 1713 517
rect 1822 485 2284 525
rect 2442 665 2488 724
rect 2442 513 2488 525
rect 1667 439 1713 471
rect 1320 405 1588 425
rect 1320 359 1335 405
rect 1569 359 1588 405
rect 1667 393 1731 439
rect 1777 393 1933 439
rect 1979 393 1990 439
rect 1667 392 1990 393
rect 1320 346 1588 359
rect 1320 312 1366 346
rect 752 244 848 269
rect 987 265 1366 312
rect 1667 273 1744 319
rect 1790 273 1968 319
rect 2014 273 2025 319
rect 987 244 1033 265
rect 752 198 765 244
rect 811 198 848 244
rect 903 198 914 244
rect 960 198 1033 244
rect 1667 219 1713 273
rect 2146 220 2222 485
rect 497 166 641 177
rect 49 134 95 146
rect 273 139 319 152
rect 543 152 641 166
rect 1079 173 1432 219
rect 1478 173 1713 219
rect 1880 200 2374 220
rect 1079 152 1125 173
rect 543 120 1125 152
rect 1926 173 2328 200
rect 1880 143 1926 154
rect 2328 142 2374 154
rect 2552 200 2598 212
rect 497 106 1125 120
rect 273 60 319 93
rect 1197 81 1208 127
rect 1254 81 1265 127
rect 1197 60 1265 81
rect 1645 81 1656 127
rect 1702 81 1713 127
rect 1645 60 1713 81
rect 2093 81 2104 127
rect 2150 81 2161 127
rect 2093 60 2161 81
rect 2552 60 2598 154
rect 0 -60 2688 60
<< labels >>
flabel metal1 s 0 724 2688 844 0 FreeSans 400 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 2552 152 2598 212 0 FreeSans 400 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel metal1 s 2238 532 2284 676 0 FreeSans 400 0 0 0 ZN
port 3 nsew default output
flabel metal1 s 74 352 324 430 0 FreeSans 400 0 0 0 EN
port 1 nsew default input
flabel metal1 s 895 358 1214 427 0 FreeSans 400 0 0 0 I
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 1822 532 1882 676 1 ZN
port 3 nsew default output
rlabel metal1 s 1822 485 2284 532 1 ZN
port 3 nsew default output
rlabel metal1 s 2146 220 2222 485 1 ZN
port 3 nsew default output
rlabel metal1 s 1880 173 2374 220 1 ZN
port 3 nsew default output
rlabel metal1 s 2328 143 2374 173 1 ZN
port 3 nsew default output
rlabel metal1 s 1880 143 1926 173 1 ZN
port 3 nsew default output
rlabel metal1 s 2328 142 2374 143 1 ZN
port 3 nsew default output
rlabel metal1 s 2442 657 2488 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2034 657 2080 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1615 657 1683 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1197 657 1265 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 291 657 359 724 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2442 604 2488 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2034 604 2080 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1615 604 1683 657 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2442 563 2488 604 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1615 563 1683 604 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2442 513 2488 563 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2552 127 2598 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 127 319 152 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2552 60 2598 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2093 60 2161 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1645 60 1713 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1197 60 1265 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 127 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2688 60 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2688 784
string GDS_END 530600
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 524022
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
