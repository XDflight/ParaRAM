magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 1206 1094
<< pwell >>
rect -86 -86 1206 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 582 573 682 939
rect 796 573 896 939
<< mvndiff >>
rect 36 294 124 333
rect 36 154 49 294
rect 95 154 124 294
rect 36 69 124 154
rect 244 294 348 333
rect 244 154 273 294
rect 319 154 348 294
rect 244 69 348 154
rect 468 294 572 333
rect 468 154 497 294
rect 543 154 572 294
rect 468 69 572 154
rect 692 285 796 333
rect 692 239 721 285
rect 767 239 796 285
rect 692 69 796 239
rect 916 294 1004 333
rect 916 154 945 294
rect 991 154 1004 294
rect 916 69 1004 154
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 861 582 939
rect 458 721 507 861
rect 553 721 582 861
rect 458 573 582 721
rect 682 573 796 939
rect 896 861 984 939
rect 896 721 925 861
rect 971 721 984 861
rect 896 573 984 721
<< mvndiffc >>
rect 49 154 95 294
rect 273 154 319 294
rect 497 154 543 294
rect 721 239 767 285
rect 945 154 991 294
<< mvpdiffc >>
rect 69 721 115 861
rect 507 721 553 861
rect 925 721 971 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 582 939 682 983
rect 796 939 896 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 377 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 377 458 454
rect 582 500 682 573
rect 582 454 595 500
rect 641 454 682 500
rect 582 377 682 454
rect 796 500 896 573
rect 796 454 814 500
rect 860 454 896 500
rect 796 377 896 454
rect 124 333 244 377
rect 348 333 468 377
rect 572 333 692 377
rect 796 333 916 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 595 454 641 500
rect 814 454 860 500
<< metal1 >>
rect 0 918 1120 1098
rect 69 861 115 918
rect 69 710 115 721
rect 507 861 553 872
rect 142 500 203 654
rect 507 603 553 721
rect 925 861 971 918
rect 925 710 971 721
rect 507 557 767 603
rect 142 454 157 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 590 500 642 511
rect 590 454 595 500
rect 641 454 642 500
rect 142 443 203 454
rect 49 351 543 397
rect 590 354 642 454
rect 49 294 95 351
rect 49 143 95 154
rect 273 294 319 305
rect 273 90 319 154
rect 497 294 543 351
rect 702 285 767 557
rect 814 500 866 511
rect 860 454 866 500
rect 814 354 866 454
rect 702 239 721 285
rect 702 228 767 239
rect 945 294 991 305
rect 543 154 945 182
rect 497 136 991 154
rect 0 -90 1120 90
<< labels >>
flabel metal1 s 590 354 642 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 814 354 866 511 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 B1
port 3 nsew default input
flabel metal1 s 142 443 203 654 0 FreeSans 200 0 0 0 B2
port 4 nsew default input
flabel metal1 s 0 918 1120 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 273 90 319 305 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 507 603 553 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 507 557 767 603 1 ZN
port 5 nsew default output
rlabel metal1 s 702 228 767 557 1 ZN
port 5 nsew default output
rlabel metal1 s 925 710 971 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 69 710 115 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 -90 1120 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1120 1008
string GDS_END 129106
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 125490
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
