magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -1273 113 1273 118
rect -1273 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1273 113
rect -1273 47 1273 85
rect -1273 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1273 47
rect -1273 -19 1273 19
rect -1273 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1273 -19
rect -1273 -85 1273 -47
rect -1273 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1273 -85
rect -1273 -118 1273 -113
<< via2 >>
rect -1268 85 -1240 113
rect -1202 85 -1174 113
rect -1136 85 -1108 113
rect -1070 85 -1042 113
rect -1004 85 -976 113
rect -938 85 -910 113
rect -872 85 -844 113
rect -806 85 -778 113
rect -740 85 -712 113
rect -674 85 -646 113
rect -608 85 -580 113
rect -542 85 -514 113
rect -476 85 -448 113
rect -410 85 -382 113
rect -344 85 -316 113
rect -278 85 -250 113
rect -212 85 -184 113
rect -146 85 -118 113
rect -80 85 -52 113
rect -14 85 14 113
rect 52 85 80 113
rect 118 85 146 113
rect 184 85 212 113
rect 250 85 278 113
rect 316 85 344 113
rect 382 85 410 113
rect 448 85 476 113
rect 514 85 542 113
rect 580 85 608 113
rect 646 85 674 113
rect 712 85 740 113
rect 778 85 806 113
rect 844 85 872 113
rect 910 85 938 113
rect 976 85 1004 113
rect 1042 85 1070 113
rect 1108 85 1136 113
rect 1174 85 1202 113
rect 1240 85 1268 113
rect -1268 19 -1240 47
rect -1202 19 -1174 47
rect -1136 19 -1108 47
rect -1070 19 -1042 47
rect -1004 19 -976 47
rect -938 19 -910 47
rect -872 19 -844 47
rect -806 19 -778 47
rect -740 19 -712 47
rect -674 19 -646 47
rect -608 19 -580 47
rect -542 19 -514 47
rect -476 19 -448 47
rect -410 19 -382 47
rect -344 19 -316 47
rect -278 19 -250 47
rect -212 19 -184 47
rect -146 19 -118 47
rect -80 19 -52 47
rect -14 19 14 47
rect 52 19 80 47
rect 118 19 146 47
rect 184 19 212 47
rect 250 19 278 47
rect 316 19 344 47
rect 382 19 410 47
rect 448 19 476 47
rect 514 19 542 47
rect 580 19 608 47
rect 646 19 674 47
rect 712 19 740 47
rect 778 19 806 47
rect 844 19 872 47
rect 910 19 938 47
rect 976 19 1004 47
rect 1042 19 1070 47
rect 1108 19 1136 47
rect 1174 19 1202 47
rect 1240 19 1268 47
rect -1268 -47 -1240 -19
rect -1202 -47 -1174 -19
rect -1136 -47 -1108 -19
rect -1070 -47 -1042 -19
rect -1004 -47 -976 -19
rect -938 -47 -910 -19
rect -872 -47 -844 -19
rect -806 -47 -778 -19
rect -740 -47 -712 -19
rect -674 -47 -646 -19
rect -608 -47 -580 -19
rect -542 -47 -514 -19
rect -476 -47 -448 -19
rect -410 -47 -382 -19
rect -344 -47 -316 -19
rect -278 -47 -250 -19
rect -212 -47 -184 -19
rect -146 -47 -118 -19
rect -80 -47 -52 -19
rect -14 -47 14 -19
rect 52 -47 80 -19
rect 118 -47 146 -19
rect 184 -47 212 -19
rect 250 -47 278 -19
rect 316 -47 344 -19
rect 382 -47 410 -19
rect 448 -47 476 -19
rect 514 -47 542 -19
rect 580 -47 608 -19
rect 646 -47 674 -19
rect 712 -47 740 -19
rect 778 -47 806 -19
rect 844 -47 872 -19
rect 910 -47 938 -19
rect 976 -47 1004 -19
rect 1042 -47 1070 -19
rect 1108 -47 1136 -19
rect 1174 -47 1202 -19
rect 1240 -47 1268 -19
rect -1268 -113 -1240 -85
rect -1202 -113 -1174 -85
rect -1136 -113 -1108 -85
rect -1070 -113 -1042 -85
rect -1004 -113 -976 -85
rect -938 -113 -910 -85
rect -872 -113 -844 -85
rect -806 -113 -778 -85
rect -740 -113 -712 -85
rect -674 -113 -646 -85
rect -608 -113 -580 -85
rect -542 -113 -514 -85
rect -476 -113 -448 -85
rect -410 -113 -382 -85
rect -344 -113 -316 -85
rect -278 -113 -250 -85
rect -212 -113 -184 -85
rect -146 -113 -118 -85
rect -80 -113 -52 -85
rect -14 -113 14 -85
rect 52 -113 80 -85
rect 118 -113 146 -85
rect 184 -113 212 -85
rect 250 -113 278 -85
rect 316 -113 344 -85
rect 382 -113 410 -85
rect 448 -113 476 -85
rect 514 -113 542 -85
rect 580 -113 608 -85
rect 646 -113 674 -85
rect 712 -113 740 -85
rect 778 -113 806 -85
rect 844 -113 872 -85
rect 910 -113 938 -85
rect 976 -113 1004 -85
rect 1042 -113 1070 -85
rect 1108 -113 1136 -85
rect 1174 -113 1202 -85
rect 1240 -113 1268 -85
<< metal3 >>
rect -1273 113 1273 118
rect -1273 85 -1268 113
rect -1240 85 -1202 113
rect -1174 85 -1136 113
rect -1108 85 -1070 113
rect -1042 85 -1004 113
rect -976 85 -938 113
rect -910 85 -872 113
rect -844 85 -806 113
rect -778 85 -740 113
rect -712 85 -674 113
rect -646 85 -608 113
rect -580 85 -542 113
rect -514 85 -476 113
rect -448 85 -410 113
rect -382 85 -344 113
rect -316 85 -278 113
rect -250 85 -212 113
rect -184 85 -146 113
rect -118 85 -80 113
rect -52 85 -14 113
rect 14 85 52 113
rect 80 85 118 113
rect 146 85 184 113
rect 212 85 250 113
rect 278 85 316 113
rect 344 85 382 113
rect 410 85 448 113
rect 476 85 514 113
rect 542 85 580 113
rect 608 85 646 113
rect 674 85 712 113
rect 740 85 778 113
rect 806 85 844 113
rect 872 85 910 113
rect 938 85 976 113
rect 1004 85 1042 113
rect 1070 85 1108 113
rect 1136 85 1174 113
rect 1202 85 1240 113
rect 1268 85 1273 113
rect -1273 47 1273 85
rect -1273 19 -1268 47
rect -1240 19 -1202 47
rect -1174 19 -1136 47
rect -1108 19 -1070 47
rect -1042 19 -1004 47
rect -976 19 -938 47
rect -910 19 -872 47
rect -844 19 -806 47
rect -778 19 -740 47
rect -712 19 -674 47
rect -646 19 -608 47
rect -580 19 -542 47
rect -514 19 -476 47
rect -448 19 -410 47
rect -382 19 -344 47
rect -316 19 -278 47
rect -250 19 -212 47
rect -184 19 -146 47
rect -118 19 -80 47
rect -52 19 -14 47
rect 14 19 52 47
rect 80 19 118 47
rect 146 19 184 47
rect 212 19 250 47
rect 278 19 316 47
rect 344 19 382 47
rect 410 19 448 47
rect 476 19 514 47
rect 542 19 580 47
rect 608 19 646 47
rect 674 19 712 47
rect 740 19 778 47
rect 806 19 844 47
rect 872 19 910 47
rect 938 19 976 47
rect 1004 19 1042 47
rect 1070 19 1108 47
rect 1136 19 1174 47
rect 1202 19 1240 47
rect 1268 19 1273 47
rect -1273 -19 1273 19
rect -1273 -47 -1268 -19
rect -1240 -47 -1202 -19
rect -1174 -47 -1136 -19
rect -1108 -47 -1070 -19
rect -1042 -47 -1004 -19
rect -976 -47 -938 -19
rect -910 -47 -872 -19
rect -844 -47 -806 -19
rect -778 -47 -740 -19
rect -712 -47 -674 -19
rect -646 -47 -608 -19
rect -580 -47 -542 -19
rect -514 -47 -476 -19
rect -448 -47 -410 -19
rect -382 -47 -344 -19
rect -316 -47 -278 -19
rect -250 -47 -212 -19
rect -184 -47 -146 -19
rect -118 -47 -80 -19
rect -52 -47 -14 -19
rect 14 -47 52 -19
rect 80 -47 118 -19
rect 146 -47 184 -19
rect 212 -47 250 -19
rect 278 -47 316 -19
rect 344 -47 382 -19
rect 410 -47 448 -19
rect 476 -47 514 -19
rect 542 -47 580 -19
rect 608 -47 646 -19
rect 674 -47 712 -19
rect 740 -47 778 -19
rect 806 -47 844 -19
rect 872 -47 910 -19
rect 938 -47 976 -19
rect 1004 -47 1042 -19
rect 1070 -47 1108 -19
rect 1136 -47 1174 -19
rect 1202 -47 1240 -19
rect 1268 -47 1273 -19
rect -1273 -85 1273 -47
rect -1273 -113 -1268 -85
rect -1240 -113 -1202 -85
rect -1174 -113 -1136 -85
rect -1108 -113 -1070 -85
rect -1042 -113 -1004 -85
rect -976 -113 -938 -85
rect -910 -113 -872 -85
rect -844 -113 -806 -85
rect -778 -113 -740 -85
rect -712 -113 -674 -85
rect -646 -113 -608 -85
rect -580 -113 -542 -85
rect -514 -113 -476 -85
rect -448 -113 -410 -85
rect -382 -113 -344 -85
rect -316 -113 -278 -85
rect -250 -113 -212 -85
rect -184 -113 -146 -85
rect -118 -113 -80 -85
rect -52 -113 -14 -85
rect 14 -113 52 -85
rect 80 -113 118 -85
rect 146 -113 184 -85
rect 212 -113 250 -85
rect 278 -113 316 -85
rect 344 -113 382 -85
rect 410 -113 448 -85
rect 476 -113 514 -85
rect 542 -113 580 -85
rect 608 -113 646 -85
rect 674 -113 712 -85
rect 740 -113 778 -85
rect 806 -113 844 -85
rect 872 -113 910 -85
rect 938 -113 976 -85
rect 1004 -113 1042 -85
rect 1070 -113 1108 -85
rect 1136 -113 1174 -85
rect 1202 -113 1240 -85
rect 1268 -113 1273 -85
rect -1273 -118 1273 -113
<< properties >>
string GDS_END 1026032
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1015916
<< end >>
