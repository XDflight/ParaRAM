magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 5420 26945 5530 27585
rect 6971 26980 7314 27448
rect 12777 26945 12875 27585
rect 14274 26980 14676 27448
rect 24877 26980 26150 27562
rect 3471 21403 3477 24683
rect 9008 22243 9090 24719
rect 10845 21403 10858 24683
rect 23104 21791 23181 24052
rect 5489 18378 8806 19567
rect 12868 18378 16185 19567
rect 20706 8070 21480 8586
rect 20739 6709 20904 6756
rect 24661 5866 24705 10029
rect 25867 5253 25991 10029
rect 27119 5388 27222 10029
rect 8352 721 8594 1303
<< mvnsubdiff >>
rect 24959 27384 25043 27403
rect 24959 27244 24978 27384
rect 25024 27244 25043 27384
rect 24959 27225 25043 27244
rect 25989 27328 26073 27347
rect 25989 27188 26008 27328
rect 26054 27188 26073 27328
rect 25989 27169 26073 27188
<< mvnsubdiffcont >>
rect 24978 27244 25024 27384
rect 26008 27188 26054 27328
<< metal1 >>
rect 403 28996 537 29037
rect 403 28944 444 28996
rect 496 28944 537 28996
rect 403 28778 537 28944
rect 1634 28939 1815 29007
rect 29520 28996 29654 29037
rect 29520 28944 29561 28996
rect 29613 28944 29654 28996
rect 403 28726 444 28778
rect 496 28726 537 28778
rect 403 1155 537 28726
rect 29520 28778 29654 28944
rect 29520 28726 29561 28778
rect 29613 28726 29654 28778
rect 24967 27384 25035 27395
rect 24967 27244 24978 27384
rect 25024 27244 25035 27384
rect 24967 27233 25035 27244
rect 25997 27328 26065 27339
rect 25997 27188 26008 27328
rect 26054 27188 26065 27328
rect 25997 27177 26065 27188
rect 6826 17625 6956 17826
rect 765 17491 6956 17625
rect 765 10724 894 17491
rect 8530 17398 8660 17813
rect 1007 17264 8660 17398
rect 1007 11101 1136 17264
rect 14218 17171 14347 17797
rect 1248 17038 14347 17171
rect 15909 17248 16038 17874
rect 24704 17475 24833 17890
rect 26395 17702 26524 17904
rect 28070 17795 28861 17928
rect 26395 17568 28619 17702
rect 24704 17342 28378 17475
rect 15909 17115 28136 17248
rect 1248 11393 1377 17038
rect 1248 11266 1843 11393
rect 1007 10945 1602 11101
rect 765 10571 1360 10724
rect 1231 1158 1360 10571
rect 1473 1158 1602 10945
rect 408 1117 532 1155
rect 408 1065 444 1117
rect 496 1065 532 1117
rect 408 899 532 1065
rect 408 847 444 899
rect 496 847 532 899
rect 408 807 532 847
rect 1231 1117 1361 1158
rect 1231 1065 1270 1117
rect 1322 1065 1361 1117
rect 1231 899 1361 1065
rect 1231 847 1270 899
rect 1322 847 1361 899
rect 1231 807 1361 847
rect 1472 1117 1602 1158
rect 1472 1065 1511 1117
rect 1563 1065 1602 1117
rect 1472 899 1602 1065
rect 1472 847 1511 899
rect 1563 847 1602 899
rect 1472 807 1602 847
rect 1231 806 1360 807
rect 1473 806 1602 807
rect 1714 1158 1843 11266
rect 21015 9604 21061 9788
rect 21463 9604 21509 9789
rect 21911 9604 21957 9796
rect 21015 9558 21957 9604
rect 20764 1590 22476 1636
rect 1714 1117 1844 1158
rect 1714 1065 1753 1117
rect 1805 1065 1844 1117
rect 1714 899 1844 1065
rect 1714 847 1753 899
rect 1805 847 1844 899
rect 1714 807 1844 847
rect 1714 806 1843 807
rect 22430 439 22476 1590
rect 28007 1130 28136 17115
rect 28007 1078 28045 1130
rect 28097 1078 28136 1130
rect 28007 912 28136 1078
rect 28007 860 28045 912
rect 28097 860 28136 912
rect 28007 694 28136 860
rect 28007 642 28045 694
rect 28097 642 28136 694
rect 28007 602 28136 642
rect 28248 1130 28378 17342
rect 28248 1078 28287 1130
rect 28339 1078 28378 1130
rect 28248 912 28378 1078
rect 28248 860 28287 912
rect 28339 860 28378 912
rect 28248 694 28378 860
rect 28248 642 28287 694
rect 28339 642 28378 694
rect 28248 602 28378 642
rect 28490 1130 28619 17568
rect 28490 1078 28529 1130
rect 28581 1078 28619 1130
rect 28490 912 28619 1078
rect 28490 860 28529 912
rect 28581 860 28619 912
rect 28490 694 28619 860
rect 28490 642 28529 694
rect 28581 642 28619 694
rect 28490 602 28619 642
rect 28731 1130 28861 17795
rect 29520 1155 29654 28726
rect 28731 1078 28770 1130
rect 28822 1078 28861 1130
rect 28731 912 28861 1078
rect 28731 860 28770 912
rect 28822 860 28861 912
rect 28731 694 28861 860
rect 29525 1117 29649 1155
rect 29525 1065 29561 1117
rect 29613 1065 29649 1117
rect 29525 899 29649 1065
rect 29525 847 29561 899
rect 29613 847 29649 899
rect 29525 807 29649 847
rect 28731 642 28770 694
rect 28822 642 28861 694
rect 28731 602 28861 642
rect 403 289 9220 330
rect 403 237 8918 289
rect 8970 237 9130 289
rect 9182 237 9220 289
rect 403 185 733 237
rect 785 185 945 237
rect 997 185 9220 237
rect 27841 237 29415 330
rect 403 71 9220 185
rect 13144 144 14721 190
rect 27841 185 29059 237
rect 29111 185 29271 237
rect 29323 185 29415 237
rect 403 19 8918 71
rect 8970 19 9130 71
rect 9182 19 9220 71
rect 403 -33 733 19
rect 785 -33 945 19
rect 997 -33 9220 19
rect 403 -126 9220 -33
rect 27841 19 29415 185
rect 27841 -33 29059 19
rect 29111 -33 29271 19
rect 29323 -33 29415 19
rect 27841 -126 29415 -33
<< via1 >>
rect 444 28944 496 28996
rect 29561 28944 29613 28996
rect 444 28726 496 28778
rect 29561 28726 29613 28778
rect 444 1065 496 1117
rect 444 847 496 899
rect 1270 1065 1322 1117
rect 1270 847 1322 899
rect 1511 1065 1563 1117
rect 1511 847 1563 899
rect 1753 1065 1805 1117
rect 1753 847 1805 899
rect 28045 1078 28097 1130
rect 28045 860 28097 912
rect 28045 642 28097 694
rect 28287 1078 28339 1130
rect 28287 860 28339 912
rect 28287 642 28339 694
rect 28529 1078 28581 1130
rect 28529 860 28581 912
rect 28529 642 28581 694
rect 28770 1078 28822 1130
rect 28770 860 28822 912
rect 29561 1065 29613 1117
rect 29561 847 29613 899
rect 28770 642 28822 694
rect 8918 237 8970 289
rect 9130 237 9182 289
rect 733 185 785 237
rect 945 185 997 237
rect 29059 185 29111 237
rect 29271 185 29323 237
rect 8918 19 8970 71
rect 9130 19 9182 71
rect 733 -33 785 19
rect 945 -33 997 19
rect 29059 -33 29111 19
rect 29271 -33 29323 19
<< metal2 >>
rect 407 28998 532 29037
rect 407 28942 442 28998
rect 498 28942 532 28998
rect 407 28780 532 28942
rect 407 28724 442 28780
rect 498 28724 532 28780
rect 407 28686 532 28724
rect 645 1382 1525 30125
rect 17156 28865 17286 28998
rect 17508 28865 17637 28998
rect 18790 28865 18920 28998
rect 19146 28865 19275 28998
rect 20426 28865 20556 28998
rect 20769 28865 20898 28998
rect 22056 28865 22185 28998
rect 22416 28865 22545 28998
rect 2336 28638 2465 28772
rect 2691 28638 2821 28772
rect 4125 28638 4255 28772
rect 4488 28638 4617 28772
rect 9714 28638 9843 28772
rect 10070 28638 10199 28772
rect 11504 28638 11633 28772
rect 11866 28638 11996 28772
rect 8963 1749 9092 1966
rect 8133 1615 9092 1749
rect 403 1117 537 1157
rect 403 1065 444 1117
rect 496 1065 537 1117
rect 403 899 537 1065
rect 403 847 444 899
rect 496 847 537 899
rect 403 -1293 537 847
rect 645 237 1086 1382
rect 645 185 733 237
rect 785 185 945 237
rect 997 185 1086 237
rect 645 19 1086 185
rect 645 -33 733 19
rect 785 -33 945 19
rect 997 -33 1086 19
rect 645 -126 1086 -33
rect 1231 1117 1361 1158
rect 1231 1065 1270 1117
rect 1322 1065 1361 1117
rect 1231 899 1361 1065
rect 1231 847 1270 899
rect 1322 847 1361 899
rect 1231 807 1361 847
rect 1472 1117 1602 1158
rect 1472 1065 1511 1117
rect 1563 1065 1602 1117
rect 1472 899 1602 1065
rect 1472 847 1511 899
rect 1563 847 1602 899
rect 1472 807 1602 847
rect 300 -1332 640 -1293
rect 300 -1388 336 -1332
rect 392 -1388 548 -1332
rect 604 -1388 640 -1332
rect 300 -1426 640 -1388
rect 403 -1427 537 -1426
rect 1231 -1427 1360 807
rect 1473 -1427 1602 807
rect 1714 1117 1844 1158
rect 1714 1065 1753 1117
rect 1805 1065 1844 1117
rect 1714 899 1844 1065
rect 1714 847 1753 899
rect 1805 847 1844 899
rect 1714 807 1844 847
rect 1714 -1427 1843 807
rect 3370 -1427 3504 1518
rect 5061 -1427 5195 1518
rect 6754 -1427 6888 1518
rect 8133 -1293 8262 1615
rect 16247 1595 16375 1651
rect 8880 289 9220 1463
rect 8880 237 8918 289
rect 8970 237 9130 289
rect 9182 237 9220 289
rect 8880 71 9220 237
rect 8880 19 8918 71
rect 8970 19 9130 71
rect 9182 19 9220 71
rect 8880 -21 9220 19
rect 8028 -1332 8368 -1293
rect 8028 -1388 8064 -1332
rect 8120 -1388 8276 -1332
rect 8332 -1388 8368 -1332
rect 8028 -1426 8368 -1388
rect 8133 -1427 8262 -1426
rect 16319 -1833 16375 1595
rect 21612 -548 21965 3456
rect 28532 1382 29412 30125
rect 29525 28998 29650 29037
rect 29525 28942 29559 28998
rect 29615 28942 29650 28998
rect 29525 28780 29650 28942
rect 29525 28724 29559 28780
rect 29615 28724 29650 28780
rect 29525 28686 29650 28724
rect 28007 1130 28136 1171
rect 28007 1078 28045 1130
rect 28097 1078 28136 1130
rect 28007 912 28136 1078
rect 28007 860 28045 912
rect 28097 860 28136 912
rect 28007 694 28136 860
rect 28007 642 28045 694
rect 28097 642 28136 694
rect 22855 -1427 22989 618
rect 28007 -1427 28136 642
rect 28248 1130 28378 1171
rect 28248 1078 28287 1130
rect 28339 1078 28378 1130
rect 28248 912 28378 1078
rect 28248 860 28287 912
rect 28339 860 28378 912
rect 28248 694 28378 860
rect 28248 642 28287 694
rect 28339 642 28378 694
rect 28248 -1427 28378 642
rect 28490 1130 28619 1171
rect 28490 1078 28529 1130
rect 28581 1078 28619 1130
rect 28490 912 28619 1078
rect 28490 860 28529 912
rect 28581 860 28619 912
rect 28490 694 28619 860
rect 28490 642 28529 694
rect 28581 642 28619 694
rect 28490 -1427 28619 642
rect 28731 1130 28861 1171
rect 28731 1078 28770 1130
rect 28822 1078 28861 1130
rect 28731 912 28861 1078
rect 28731 860 28770 912
rect 28822 860 28861 912
rect 28731 694 28861 860
rect 28731 642 28770 694
rect 28822 642 28861 694
rect 28731 -1427 28861 642
rect 28971 237 29412 1382
rect 28971 185 29059 237
rect 29111 185 29271 237
rect 29323 185 29412 237
rect 28971 19 29412 185
rect 28971 -33 29059 19
rect 29111 -33 29271 19
rect 29323 -33 29412 19
rect 28971 -126 29412 -33
rect 29520 1117 29654 1157
rect 29520 1065 29561 1117
rect 29613 1065 29654 1117
rect 29520 899 29654 1065
rect 29520 847 29561 899
rect 29613 847 29654 899
rect 29520 -1293 29654 847
rect 29417 -1332 29757 -1293
rect 29417 -1388 29453 -1332
rect 29509 -1388 29665 -1332
rect 29721 -1388 29757 -1332
rect 29417 -1426 29757 -1388
rect 29520 -1427 29654 -1426
<< via2 >>
rect 442 28996 498 28998
rect 442 28944 444 28996
rect 444 28944 496 28996
rect 496 28944 498 28996
rect 442 28942 498 28944
rect 442 28778 498 28780
rect 442 28726 444 28778
rect 444 28726 496 28778
rect 496 28726 498 28778
rect 442 28724 498 28726
rect 336 -1388 392 -1332
rect 548 -1388 604 -1332
rect 8064 -1388 8120 -1332
rect 8276 -1388 8332 -1332
rect 29559 28996 29615 28998
rect 29559 28944 29561 28996
rect 29561 28944 29613 28996
rect 29613 28944 29615 28996
rect 29559 28942 29615 28944
rect 29559 28778 29615 28780
rect 29559 28726 29561 28778
rect 29561 28726 29613 28778
rect 29613 28726 29615 28778
rect 29559 28724 29615 28726
rect 29453 -1388 29509 -1332
rect 29665 -1388 29721 -1332
<< metal3 >>
rect 645 29216 29412 30125
rect 403 28998 29654 29037
rect 403 28942 442 28998
rect 498 28942 29559 28998
rect 29615 28942 29654 28998
rect 403 28780 29654 28942
rect 403 28724 442 28780
rect 498 28724 29559 28780
rect 29615 28724 29654 28780
rect 403 28686 29654 28724
rect 407 28685 533 28686
rect 29524 28685 29650 28686
rect 28110 14839 28239 14972
rect 28110 14499 28239 14632
rect 28110 14159 28239 14292
rect 28110 13819 28239 13952
rect 28110 13479 28239 13612
rect 28110 13139 28239 13272
rect 28110 12798 28239 12932
rect 28110 12458 28239 12592
rect 13919 6986 14239 7863
rect 16097 1580 16589 1668
rect 300 -1332 640 -1293
rect 300 -1388 336 -1332
rect 392 -1388 548 -1332
rect 604 -1388 640 -1332
rect 300 -1426 640 -1388
rect 8028 -1332 8368 -1293
rect 8028 -1388 8064 -1332
rect 8120 -1388 8276 -1332
rect 8332 -1388 8368 -1332
rect 8028 -1426 8368 -1388
rect 29417 -1332 29757 -1293
rect 29417 -1388 29453 -1332
rect 29509 -1388 29665 -1332
rect 29721 -1388 29757 -1332
rect 29417 -1426 29757 -1388
use M1_NACTIVE4310590548746_128x8m81  M1_NACTIVE4310590548746_128x8m81_0
timestamp 1666464484
transform 0 -1 26031 1 0 27258
box 0 0 1 1
use M1_NACTIVE4310590548746_128x8m81  M1_NACTIVE4310590548746_128x8m81_1
timestamp 1666464484
transform 0 -1 25001 1 0 27314
box 0 0 1 1
use M1_PACTIVE4310590548747_128x8m81  M1_PACTIVE4310590548747_128x8m81_0
timestamp 1666464484
transform 1 0 3487 0 1 28973
box -1734 -42 1734 42
use M1_PACTIVE4310590548747_128x8m81  M1_PACTIVE4310590548747_128x8m81_1
timestamp 1666464484
transform 1 0 10847 0 1 28973
box -1734 -42 1734 42
use M1_PACTIVE4310590548748_128x8m81  M1_PACTIVE4310590548748_128x8m81_0
timestamp 1666464484
transform 1 0 23865 0 1 28384
box -653 -42 653 42
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_0
timestamp 1666464484
transform -1 0 29587 0 1 28861
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_1
timestamp 1666464484
transform -1 0 29587 0 1 982
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_2
timestamp 1666464484
transform 1 0 470 0 1 28861
box 0 0 1 1
use M2_M1$$43375660_128x8m81  M2_M1$$43375660_128x8m81_3
timestamp 1666464484
transform 1 0 470 0 1 982
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_0
timestamp 1666464484
transform 1 0 865 0 1 102
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_1
timestamp 1666464484
transform 1 0 29191 0 1 102
box 0 0 1 1
use M2_M1$$199746604_128x8m81  M2_M1$$199746604_128x8m81_2
timestamp 1666464484
transform 1 0 9050 0 1 154
box 0 0 1 1
use M2_M1$$201262124_128x8m81  M2_M1$$201262124_128x8m81_0
timestamp 1666464484
transform 1 0 9050 0 1 263
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_0
timestamp 1666464484
transform 1 0 28796 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_1
timestamp 1666464484
transform 1 0 28555 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_2
timestamp 1666464484
transform 1 0 28313 0 1 886
box 0 0 1 1
use M2_M1$$202405932_128x8m81  M2_M1$$202405932_128x8m81_3
timestamp 1666464484
transform 1 0 28071 0 1 886
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_0
timestamp 1666464484
transform 1 0 1779 0 1 982
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_1
timestamp 1666464484
transform 1 0 1537 0 1 982
box 0 0 1 1
use M2_M1$$202406956_128x8m81  M2_M1$$202406956_128x8m81_2
timestamp 1666464484
transform 1 0 1296 0 1 982
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_0
timestamp 1666464484
transform -1 0 29587 0 1 28861
box 0 0 1 1
use M3_M2$$43368492_128x8m81_0  M3_M2$$43368492_128x8m81_0_1
timestamp 1666464484
transform 1 0 470 0 1 28861
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_0
timestamp 1666464484
transform -1 0 29587 0 1 -1360
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_1
timestamp 1666464484
transform 1 0 470 0 1 -1360
box 0 0 1 1
use M3_M2$$201255980_128x8m81  M3_M2$$201255980_128x8m81_2
timestamp 1666464484
transform 1 0 8198 0 1 -1360
box 0 0 1 1
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_0
timestamp 1666464484
transform 1 0 28972 0 1 29671
box -381 -393 381 393
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_1
timestamp 1666464484
transform 1 0 1085 0 1 29671
box -381 -393 381 393
use M3_M2$$201401388_128x8m81  M3_M2$$201401388_128x8m81_2
timestamp 1666464484
transform 1 0 28972 0 1 9689
box -381 -393 381 393
use M3_M24310590548749_128x8m81  M3_M24310590548749_128x8m81_0
timestamp 1666464484
transform 1 0 21792 0 1 -321
box -142 -142 142 142
use M3_M24310590548749_128x8m81  M3_M24310590548749_128x8m81_1
timestamp 1666464484
transform 1 0 21792 0 1 747
box -142 -142 142 142
use gen_512x8_128x8m81  gen_512x8_128x8m81_0
timestamp 1666464484
transform 1 0 14166 0 1 714
box -17790 -2370 17624 16428
use prexdec_top_128x8m81  prexdec_top_128x8m81_0
timestamp 1666464484
transform 1 0 1357 0 1 17581
box 36 -1 27315 12544
use ypredec1_128x8m81  ypredec1_128x8m81_0
timestamp 1666464484
transform 1 0 1561 0 1 560
box 179 76 26678 16532
<< labels >>
flabel metal3 s 8281 -1000 8281 -1000 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 8281 -352 8281 -352 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
rlabel metal3 s 28175 14906 28175 14906 4 RYS[7]
port 3 nsew
rlabel metal3 s 28175 14565 28175 14565 4 RYS[6]
port 4 nsew
rlabel metal3 s 28175 14225 28175 14225 4 RYS[5]
port 5 nsew
rlabel metal3 s 28175 13885 28175 13885 4 RYS[4]
port 6 nsew
rlabel metal3 s 28175 13545 28175 13545 4 RYS[3]
port 7 nsew
rlabel metal3 s 28175 13205 28175 13205 4 RYS[2]
port 8 nsew
rlabel metal3 s 28175 12865 28175 12865 4 RYS[1]
port 9 nsew
rlabel metal3 s 28175 12525 28175 12525 4 RYS[0]
port 10 nsew
rlabel metal3 s 1805 12525 1805 12525 4 LYS[0]
port 11 nsew
rlabel metal3 s 1805 12865 1805 12865 4 LYS[1]
port 12 nsew
rlabel metal3 s 1805 13205 1805 13205 4 LYS[2]
port 13 nsew
rlabel metal3 s 1805 13545 1805 13545 4 LYS[3]
port 14 nsew
rlabel metal3 s 1805 14565 1805 14565 4 LYS[6]
port 15 nsew
rlabel metal3 s 1805 14225 1805 14225 4 LYS[5]
port 16 nsew
rlabel metal3 s 1805 13885 1805 13885 4 LYS[4]
port 17 nsew
rlabel metal3 s 26861 29671 26861 29671 4 men
port 18 nsew
rlabel metal3 s 1805 14906 1805 14906 4 LYS[7]
port 19 nsew
rlabel metal3 s 27957 5019 27957 5019 4 tblhl
port 20 nsew
flabel metal3 s 6236 9021 6236 9021 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 18161 6236 18161 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 3499 6236 3499 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 1395 6236 1395 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 8281 1059 8281 1059 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 18981 6236 18981 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 24007 6236 24007 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 2448 6236 2448 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 28103 6236 28103 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 26066 6236 26066 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal3 s 6236 6539 6236 6539 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 15970 6236 15970 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 27112 6236 27112 0 FreeSans 2000 0 0 0 VDD
port 2 nsew
flabel metal3 s 6236 20288 6236 20288 0 FreeSans 2000 0 0 0 VSS
port 1 nsew
flabel metal2 s 16356 -1340 16356 -1340 0 FreeSans 1000 0 0 0 IGWEN
port 21 nsew
rlabel metal2 s 9726 28748 9726 28748 4 xb[3]
port 22 nsew
rlabel metal2 s 10163 28755 10163 28755 4 xb[2]
port 23 nsew
rlabel metal2 s 11966 28730 11966 28730 4 xb[0]
port 24 nsew
rlabel metal2 s 17221 28931 17221 28931 4 xa[7]
port 25 nsew
rlabel metal2 s 17572 28931 17572 28931 4 xa[6]
port 26 nsew
rlabel metal2 s 18855 28931 18855 28931 4 xa[5]
port 27 nsew
rlabel metal2 s 19211 28931 19211 28931 4 xa[4]
port 28 nsew
rlabel metal2 s 20491 28931 20491 28931 4 xa[3]
port 29 nsew
rlabel metal2 s 20833 28931 20833 28931 4 xa[2]
port 30 nsew
rlabel metal2 s 6821 -1360 6821 -1360 4 A[0]
port 31 nsew
rlabel metal2 s 22924 -1360 22924 -1360 4 CEN
port 32 nsew
rlabel metal2 s 11527 28712 11527 28712 4 xb[1]
port 33 nsew
rlabel metal2 s 10135 28705 10135 28705 4 xb[2]
port 23 nsew
rlabel metal2 s 11931 28700 11931 28700 4 xb[0]
port 24 nsew
rlabel metal2 s 2400 28705 2400 28705 4 xc[3]
port 34 nsew
rlabel metal2 s 4190 28700 4190 28700 4 xc[1]
port 35 nsew
rlabel metal2 s 2756 28705 2756 28705 4 xc[2]
port 36 nsew
rlabel metal2 s 4552 28700 4552 28700 4 xc[0]
port 37 nsew
rlabel metal2 s 22480 28931 22480 28931 4 xa[0]
port 38 nsew
rlabel metal2 s 22120 28931 22120 28931 4 xa[1]
port 39 nsew
rlabel metal2 s 1296 -1360 1296 -1360 4 A[9]
port 40 nsew
rlabel metal2 s 1779 -1360 1779 -1360 4 A[7]
port 41 nsew
rlabel metal2 s 470 -1360 470 -1360 4 CLK
port 42 nsew
rlabel metal2 s 11569 28700 11569 28700 4 xb[1]
port 33 nsew
rlabel metal2 s 9779 28705 9779 28705 4 xb[3]
port 22 nsew
rlabel metal2 s 3437 -1360 3437 -1360 4 A[2]
port 43 nsew
rlabel metal2 s 5128 -1360 5128 -1360 4 A[1]
port 44 nsew
rlabel metal2 s 28071 -1360 28071 -1360 4 A[6]
port 45 nsew
rlabel metal2 s 28796 -1360 28796 -1360 4 A[3]
port 46 nsew
rlabel metal2 s 28555 -1360 28555 -1360 4 A[4]
port 47 nsew
rlabel metal2 s 28313 -1360 28313 -1360 4 A[5]
port 48 nsew
rlabel metal2 s 1537 -1360 1537 -1360 4 A[8]
port 49 nsew
flabel metal1 s 22454 1053 22454 1053 0 FreeSans 1000 0 0 0 GWE
port 50 nsew
<< properties >>
string GDS_END 2297844
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2287270
string path 80.485 8.120 82.945 8.120 
<< end >>
