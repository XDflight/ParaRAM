magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -220 -636 221 636
<< nsubdiff >>
rect -77 431 78 488
rect -77 385 -23 431
rect 23 385 78 431
rect -77 268 78 385
rect -77 222 -23 268
rect 23 222 78 268
rect -77 105 78 222
rect -77 59 -23 105
rect 23 59 78 105
rect -77 -59 78 59
rect -77 -105 -23 -59
rect 23 -105 78 -59
rect -77 -222 78 -105
rect -77 -268 -23 -222
rect 23 -268 78 -222
rect -77 -385 78 -268
rect -77 -431 -23 -385
rect 23 -431 78 -385
rect -77 -488 78 -431
<< nsubdiffcont >>
rect -23 385 23 431
rect -23 222 23 268
rect -23 59 23 105
rect -23 -105 23 -59
rect -23 -268 23 -222
rect -23 -431 23 -385
<< metal1 >>
rect -57 431 58 468
rect -57 385 -23 431
rect 23 385 58 431
rect -57 268 58 385
rect -57 222 -23 268
rect 23 222 58 268
rect -57 105 58 222
rect -57 59 -23 105
rect 23 59 58 105
rect -57 -59 58 59
rect -57 -105 -23 -59
rect 23 -105 58 -59
rect -57 -222 58 -105
rect -57 -268 -23 -222
rect 23 -268 58 -222
rect -57 -385 58 -268
rect -57 -431 -23 -385
rect 23 -431 58 -385
rect -57 -468 58 -431
<< properties >>
string GDS_END 226048
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 225404
<< end >>
