magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 982 1094
<< pwell >>
rect -86 -86 982 453
<< mvnmos >>
rect 124 69 244 227
rect 348 69 468 227
rect 572 69 692 227
<< mvpmos >>
rect 144 573 244 939
rect 358 573 458 939
rect 572 573 672 939
<< mvndiff >>
rect 36 193 124 227
rect 36 147 49 193
rect 95 147 124 193
rect 36 69 124 147
rect 244 193 348 227
rect 244 147 273 193
rect 319 147 348 193
rect 244 69 348 147
rect 468 193 572 227
rect 468 147 497 193
rect 543 147 572 193
rect 468 69 572 147
rect 692 193 780 227
rect 692 147 721 193
rect 767 147 780 193
rect 692 69 780 147
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 573 358 939
rect 458 573 572 939
rect 672 861 760 939
rect 672 721 701 861
rect 747 721 760 861
rect 672 573 760 721
<< mvndiffc >>
rect 49 147 95 193
rect 273 147 319 193
rect 497 147 543 193
rect 721 147 767 193
<< mvpdiffc >>
rect 69 721 115 861
rect 701 721 747 861
<< polysilicon >>
rect 144 939 244 983
rect 358 939 458 983
rect 572 939 672 983
rect 144 500 244 573
rect 144 454 157 500
rect 203 454 244 500
rect 144 271 244 454
rect 358 500 458 573
rect 358 454 371 500
rect 417 454 458 500
rect 358 271 458 454
rect 572 500 672 573
rect 572 454 590 500
rect 636 454 672 500
rect 572 271 672 454
rect 124 227 244 271
rect 348 227 468 271
rect 572 227 692 271
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
<< polycontact >>
rect 157 454 203 500
rect 371 454 417 500
rect 590 454 636 500
<< metal1 >>
rect 0 918 896 1098
rect 69 861 115 918
rect 69 710 115 721
rect 701 861 767 872
rect 747 721 767 861
rect 142 500 203 542
rect 142 454 157 500
rect 360 500 428 542
rect 360 454 371 500
rect 417 454 428 500
rect 590 500 642 511
rect 636 454 642 500
rect 142 443 203 454
rect 590 354 642 454
rect 701 296 767 721
rect 273 250 767 296
rect 49 193 95 204
rect 49 90 95 147
rect 273 193 319 250
rect 273 136 319 147
rect 497 193 543 204
rect 497 90 543 147
rect 721 193 767 250
rect 721 136 767 147
rect 0 -90 896 90
<< labels >>
flabel metal1 s 590 354 642 511 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 360 454 428 542 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 142 443 203 542 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 918 896 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 497 90 543 204 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 701 296 767 872 0 FreeSans 200 0 0 0 ZN
port 4 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 273 250 767 296 1 ZN
port 4 nsew default output
rlabel metal1 s 721 136 767 250 1 ZN
port 4 nsew default output
rlabel metal1 s 273 136 319 250 1 ZN
port 4 nsew default output
rlabel metal1 s 69 710 115 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 49 90 95 204 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 896 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string GDS_END 86456
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 83686
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
