magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 1448 616
<< mvpmos >>
rect 0 0 120 496
rect 224 0 344 496
rect 448 0 568 496
rect 672 0 792 496
rect 896 0 1016 496
rect 1120 0 1240 496
<< mvpdiff >>
rect -88 483 0 496
rect -88 437 -75 483
rect -29 437 0 483
rect -88 377 0 437
rect -88 331 -75 377
rect -29 331 0 377
rect -88 271 0 331
rect -88 225 -75 271
rect -29 225 0 271
rect -88 165 0 225
rect -88 119 -75 165
rect -29 119 0 165
rect -88 59 0 119
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 483 224 496
rect 120 437 149 483
rect 195 437 224 483
rect 120 377 224 437
rect 120 331 149 377
rect 195 331 224 377
rect 120 271 224 331
rect 120 225 149 271
rect 195 225 224 271
rect 120 165 224 225
rect 120 119 149 165
rect 195 119 224 165
rect 120 59 224 119
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 483 448 496
rect 344 437 373 483
rect 419 437 448 483
rect 344 377 448 437
rect 344 331 373 377
rect 419 331 448 377
rect 344 271 448 331
rect 344 225 373 271
rect 419 225 448 271
rect 344 165 448 225
rect 344 119 373 165
rect 419 119 448 165
rect 344 59 448 119
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 483 672 496
rect 568 437 597 483
rect 643 437 672 483
rect 568 377 672 437
rect 568 331 597 377
rect 643 331 672 377
rect 568 271 672 331
rect 568 225 597 271
rect 643 225 672 271
rect 568 165 672 225
rect 568 119 597 165
rect 643 119 672 165
rect 568 59 672 119
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 483 896 496
rect 792 437 821 483
rect 867 437 896 483
rect 792 377 896 437
rect 792 331 821 377
rect 867 331 896 377
rect 792 271 896 331
rect 792 225 821 271
rect 867 225 896 271
rect 792 165 896 225
rect 792 119 821 165
rect 867 119 896 165
rect 792 59 896 119
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 483 1120 496
rect 1016 437 1045 483
rect 1091 437 1120 483
rect 1016 377 1120 437
rect 1016 331 1045 377
rect 1091 331 1120 377
rect 1016 271 1120 331
rect 1016 225 1045 271
rect 1091 225 1120 271
rect 1016 165 1120 225
rect 1016 119 1045 165
rect 1091 119 1120 165
rect 1016 59 1120 119
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 483 1328 496
rect 1240 437 1269 483
rect 1315 437 1328 483
rect 1240 377 1328 437
rect 1240 331 1269 377
rect 1315 331 1328 377
rect 1240 271 1328 331
rect 1240 225 1269 271
rect 1315 225 1328 271
rect 1240 165 1328 225
rect 1240 119 1269 165
rect 1315 119 1328 165
rect 1240 59 1328 119
rect 1240 13 1269 59
rect 1315 13 1328 59
rect 1240 0 1328 13
<< mvpdiffc >>
rect -75 437 -29 483
rect -75 331 -29 377
rect -75 225 -29 271
rect -75 119 -29 165
rect -75 13 -29 59
rect 149 437 195 483
rect 149 331 195 377
rect 149 225 195 271
rect 149 119 195 165
rect 149 13 195 59
rect 373 437 419 483
rect 373 331 419 377
rect 373 225 419 271
rect 373 119 419 165
rect 373 13 419 59
rect 597 437 643 483
rect 597 331 643 377
rect 597 225 643 271
rect 597 119 643 165
rect 597 13 643 59
rect 821 437 867 483
rect 821 331 867 377
rect 821 225 867 271
rect 821 119 867 165
rect 821 13 867 59
rect 1045 437 1091 483
rect 1045 331 1091 377
rect 1045 225 1091 271
rect 1045 119 1091 165
rect 1045 13 1091 59
rect 1269 437 1315 483
rect 1269 331 1315 377
rect 1269 225 1315 271
rect 1269 119 1315 165
rect 1269 13 1315 59
<< polysilicon >>
rect 0 496 120 540
rect 224 496 344 540
rect 448 496 568 540
rect 672 496 792 540
rect 896 496 1016 540
rect 1120 496 1240 540
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
<< metal1 >>
rect -75 483 -29 496
rect -75 377 -29 437
rect -75 271 -29 331
rect -75 165 -29 225
rect -75 59 -29 119
rect -75 0 -29 13
rect 149 483 195 496
rect 149 377 195 437
rect 149 271 195 331
rect 149 165 195 225
rect 149 59 195 119
rect 149 0 195 13
rect 373 483 419 496
rect 373 377 419 437
rect 373 271 419 331
rect 373 165 419 225
rect 373 59 419 119
rect 373 0 419 13
rect 597 483 643 496
rect 597 377 643 437
rect 597 271 643 331
rect 597 165 643 225
rect 597 59 643 119
rect 597 0 643 13
rect 821 483 867 496
rect 821 377 867 437
rect 821 271 867 331
rect 821 165 867 225
rect 821 59 867 119
rect 821 0 867 13
rect 1045 483 1091 496
rect 1045 377 1091 437
rect 1045 271 1091 331
rect 1045 165 1091 225
rect 1045 59 1091 119
rect 1045 0 1091 13
rect 1269 483 1315 496
rect 1269 377 1315 437
rect 1269 271 1315 331
rect 1269 165 1315 225
rect 1269 59 1315 119
rect 1269 0 1315 13
<< labels >>
flabel metal1 s -52 248 -52 248 0 FreeSans 400 0 0 0 S
flabel metal1 s 1292 248 1292 248 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 248 172 248 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 248 396 248 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 248 620 248 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 248 844 248 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 248 1068 248 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 536344
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 531234
<< end >>
