magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 5600 844
rect 49 506 95 724
rect 477 600 523 724
rect 925 600 971 724
rect 1373 600 1419 724
rect 1821 506 1867 724
rect 2065 562 2111 676
rect 2269 608 2315 724
rect 2493 562 2539 676
rect 2717 608 2763 724
rect 2941 562 2987 676
rect 3165 608 3211 724
rect 3389 562 3435 676
rect 3613 608 3659 724
rect 3837 562 3883 676
rect 4061 608 4107 724
rect 4285 562 4331 676
rect 4509 608 4555 724
rect 4733 562 4779 676
rect 4957 608 5003 724
rect 5181 562 5227 676
rect 124 342 1637 430
rect 2065 446 5227 562
rect 5405 506 5451 724
rect 3550 302 3730 446
rect 38 60 106 153
rect 486 60 554 153
rect 934 60 1002 153
rect 1382 60 1450 153
rect 2065 186 5247 302
rect 1830 60 1898 153
rect 2065 135 2117 186
rect 2278 60 2346 140
rect 2513 135 2559 186
rect 2726 60 2794 140
rect 2961 135 3007 186
rect 3174 60 3242 140
rect 3409 135 3455 186
rect 3622 60 3690 140
rect 3857 135 3903 186
rect 4070 60 4138 140
rect 4305 135 4351 186
rect 4518 60 4586 140
rect 4753 135 4799 186
rect 4966 60 5034 140
rect 5201 135 5247 186
rect 5414 60 5482 153
rect 0 -60 5600 60
<< obsm1 >>
rect 253 552 299 676
rect 701 552 747 676
rect 1149 552 1195 676
rect 1597 552 1643 676
rect 253 506 1754 552
rect 1707 394 1754 506
rect 1707 348 3302 394
rect 1707 250 1754 348
rect 3912 348 5396 394
rect 273 203 1754 250
rect 273 135 319 203
rect 721 135 767 203
rect 1169 135 1215 203
rect 1617 135 1663 203
<< labels >>
rlabel metal1 s 124 342 1637 430 6 I
port 1 nsew default input
rlabel metal1 s 5181 562 5227 676 6 Z
port 2 nsew default output
rlabel metal1 s 4733 562 4779 676 6 Z
port 2 nsew default output
rlabel metal1 s 4285 562 4331 676 6 Z
port 2 nsew default output
rlabel metal1 s 3837 562 3883 676 6 Z
port 2 nsew default output
rlabel metal1 s 3389 562 3435 676 6 Z
port 2 nsew default output
rlabel metal1 s 2941 562 2987 676 6 Z
port 2 nsew default output
rlabel metal1 s 2493 562 2539 676 6 Z
port 2 nsew default output
rlabel metal1 s 2065 562 2111 676 6 Z
port 2 nsew default output
rlabel metal1 s 2065 446 5227 562 6 Z
port 2 nsew default output
rlabel metal1 s 3550 302 3730 446 6 Z
port 2 nsew default output
rlabel metal1 s 2065 186 5247 302 6 Z
port 2 nsew default output
rlabel metal1 s 5201 135 5247 186 6 Z
port 2 nsew default output
rlabel metal1 s 4753 135 4799 186 6 Z
port 2 nsew default output
rlabel metal1 s 4305 135 4351 186 6 Z
port 2 nsew default output
rlabel metal1 s 3857 135 3903 186 6 Z
port 2 nsew default output
rlabel metal1 s 3409 135 3455 186 6 Z
port 2 nsew default output
rlabel metal1 s 2961 135 3007 186 6 Z
port 2 nsew default output
rlabel metal1 s 2513 135 2559 186 6 Z
port 2 nsew default output
rlabel metal1 s 2065 135 2117 186 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 5600 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 608 5451 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4957 608 5003 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4509 608 4555 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 4061 608 4107 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3613 608 3659 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3165 608 3211 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2717 608 2763 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2269 608 2315 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 608 1867 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 608 1419 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 608 971 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 608 523 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 608 95 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 600 5451 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 600 1867 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1373 600 1419 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 925 600 971 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 477 600 523 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 600 95 608 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5405 506 5451 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1821 506 1867 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 49 506 95 600 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 5414 140 5482 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 140 1898 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 140 1450 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 140 1002 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 140 554 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 38 140 106 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 5414 60 5482 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4966 60 5034 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4518 60 4586 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 4070 60 4138 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3622 60 3690 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3174 60 3242 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2726 60 2794 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2278 60 2346 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1830 60 1898 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1382 60 1450 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 934 60 1002 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 140 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5600 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5600 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1345084
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1333176
<< end >>
