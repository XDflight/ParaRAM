magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 688
<< mvpmos >>
rect 0 0 120 568
rect 224 0 344 568
<< mvpdiff >>
rect -88 555 0 568
rect -88 509 -75 555
rect -29 509 0 555
rect -88 431 0 509
rect -88 385 -75 431
rect -29 385 0 431
rect -88 307 0 385
rect -88 261 -75 307
rect -29 261 0 307
rect -88 183 0 261
rect -88 137 -75 183
rect -29 137 0 183
rect -88 59 0 137
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 555 224 568
rect 120 509 149 555
rect 195 509 224 555
rect 120 431 224 509
rect 120 385 149 431
rect 195 385 224 431
rect 120 307 224 385
rect 120 261 149 307
rect 195 261 224 307
rect 120 183 224 261
rect 120 137 149 183
rect 195 137 224 183
rect 120 59 224 137
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 555 432 568
rect 344 509 373 555
rect 419 509 432 555
rect 344 431 432 509
rect 344 385 373 431
rect 419 385 432 431
rect 344 307 432 385
rect 344 261 373 307
rect 419 261 432 307
rect 344 183 432 261
rect 344 137 373 183
rect 419 137 432 183
rect 344 59 432 137
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 509 -29 555
rect -75 385 -29 431
rect -75 261 -29 307
rect -75 137 -29 183
rect -75 13 -29 59
rect 149 509 195 555
rect 149 385 195 431
rect 149 261 195 307
rect 149 137 195 183
rect 149 13 195 59
rect 373 509 419 555
rect 373 385 419 431
rect 373 261 419 307
rect 373 137 419 183
rect 373 13 419 59
<< polysilicon >>
rect 0 568 120 612
rect 224 568 344 612
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 555 -29 568
rect -75 431 -29 509
rect -75 307 -29 385
rect -75 183 -29 261
rect -75 59 -29 137
rect -75 0 -29 13
rect 149 555 195 568
rect 149 431 195 509
rect 149 307 195 385
rect 149 183 195 261
rect 149 59 195 137
rect 149 0 195 13
rect 373 555 419 568
rect 373 431 419 509
rect 373 307 419 385
rect 373 183 419 261
rect 373 59 419 137
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 284 -52 284 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 284 396 284 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 284 172 284 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 611610
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 609308
<< end >>
