magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 454 89 527
rect 193 454 313 527
rect 417 454 537 527
rect 641 454 761 527
rect 865 454 985 527
rect 1089 454 1209 527
rect 1313 454 1433 527
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 641 -74 761 -1
rect 865 -74 985 -1
rect 1089 -74 1209 -1
rect 1313 -74 1433 -1
use nmos_5p04310589983225_64x8m81  nmos_5p04310589983225_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 1552 498
<< properties >>
string GDS_END 324704
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 323686
<< end >>
