magic
tech gf180mcuC
timestamp 1667403421
<< metal1 >>
rect 0 147 260 159
rect 28 106 33 147
rect 89 106 94 147
rect 145 121 150 147
rect 52 80 75 86
rect 38 67 48 73
rect 67 47 73 80
rect 177 106 182 147
rect 110 80 131 86
rect 65 41 75 47
rect 110 46 116 80
rect 153 80 163 86
rect 209 86 214 140
rect 226 106 231 147
rect 243 100 248 140
rect 243 93 253 100
rect 243 92 252 93
rect 209 80 238 86
rect 108 40 118 46
rect 28 9 33 33
rect 89 9 94 25
rect 145 9 150 33
rect 177 9 182 26
rect 231 43 236 80
rect 209 38 236 43
rect 209 16 214 38
rect 226 9 231 33
rect 243 16 248 92
rect 0 -3 260 9
<< obsm1 >>
rect 11 49 16 140
rect 61 101 66 140
rect 117 121 122 140
rect 99 116 122 121
rect 28 96 66 101
rect 28 86 33 96
rect 81 93 91 99
rect 21 80 33 86
rect 10 39 16 49
rect 28 47 33 80
rect 83 47 89 93
rect 99 71 104 116
rect 134 93 144 99
rect 162 97 167 140
rect 98 66 104 71
rect 28 42 48 47
rect 11 16 16 39
rect 40 33 48 42
rect 81 41 91 47
rect 98 34 103 66
rect 136 73 142 93
rect 162 92 178 97
rect 172 73 178 92
rect 135 67 146 73
rect 162 68 178 73
rect 136 66 144 67
rect 121 54 131 60
rect 162 52 168 68
rect 181 60 187 62
rect 194 60 199 140
rect 179 54 189 60
rect 194 54 223 60
rect 40 28 66 33
rect 98 29 125 34
rect 61 16 66 28
rect 117 28 125 29
rect 117 16 122 28
rect 162 16 167 52
rect 181 37 187 54
rect 179 31 189 37
rect 194 16 199 54
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 58 154 66 155
rect 82 154 90 155
rect 106 154 114 155
rect 130 154 138 155
rect 154 154 162 155
rect 178 154 186 155
rect 202 154 210 155
rect 226 154 234 155
rect 9 148 19 154
rect 33 148 43 154
rect 57 148 67 154
rect 81 148 91 154
rect 105 148 115 154
rect 129 148 139 154
rect 153 148 163 154
rect 177 148 187 154
rect 201 148 211 154
rect 225 148 235 154
rect 10 147 18 148
rect 34 147 42 148
rect 58 147 66 148
rect 82 147 90 148
rect 106 147 114 148
rect 130 147 138 148
rect 154 147 162 148
rect 178 147 186 148
rect 202 147 210 148
rect 226 147 234 148
rect 244 99 252 100
rect 243 93 253 99
rect 65 86 74 87
rect 121 86 131 87
rect 154 86 162 87
rect 65 80 163 86
rect 65 79 74 80
rect 121 79 131 80
rect 154 79 162 80
rect 38 73 48 74
rect 35 67 51 73
rect 38 66 48 67
rect 244 92 252 93
rect 229 86 237 87
rect 228 80 238 86
rect 229 79 237 80
rect 10 8 18 9
rect 34 8 42 9
rect 58 8 66 9
rect 82 8 90 9
rect 106 8 114 9
rect 130 8 138 9
rect 154 8 162 9
rect 178 8 186 9
rect 202 8 210 9
rect 226 8 234 9
rect 9 2 19 8
rect 33 2 43 8
rect 57 2 67 8
rect 81 2 91 8
rect 105 2 115 8
rect 129 2 139 8
rect 153 2 163 8
rect 177 2 187 8
rect 201 2 211 8
rect 225 2 235 8
rect 10 1 18 2
rect 34 1 42 2
rect 58 1 66 2
rect 82 1 90 2
rect 106 1 114 2
rect 130 1 138 2
rect 154 1 162 2
rect 178 1 186 2
rect 202 1 210 2
rect 226 1 234 2
<< obsm2 >>
rect 135 99 143 100
rect 134 93 198 99
rect 135 92 143 93
rect 136 73 144 74
rect 135 67 145 73
rect 136 66 144 67
rect 122 60 130 61
rect 161 60 169 61
rect 192 60 198 93
rect 214 60 222 61
rect 121 54 171 60
rect 192 54 223 60
rect 122 53 130 54
rect 161 53 169 54
rect 214 53 222 54
rect 9 47 17 48
rect 82 47 90 48
rect 8 41 91 47
rect 9 40 17 41
rect 82 40 90 41
rect 180 37 188 38
rect 116 34 124 35
rect 170 34 189 37
rect 115 31 189 34
rect 115 30 188 31
rect 115 28 176 30
rect 116 27 124 28
<< labels >>
rlabel metal2 s 65 79 74 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 121 79 131 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 154 79 162 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 65 80 163 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 67 41 73 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 65 41 75 47 6 CLK
port 1 nsew clock input
rlabel metal1 s 52 80 75 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 110 40 116 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 108 40 118 46 6 CLK
port 1 nsew clock input
rlabel metal1 s 110 80 131 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 153 80 163 86 6 CLK
port 1 nsew clock input
rlabel metal2 s 38 66 48 74 6 D
port 2 nsew signal input
rlabel metal2 s 35 67 51 73 6 D
port 2 nsew signal input
rlabel metal1 s 38 67 48 73 6 D
port 2 nsew signal input
rlabel metal2 s 244 92 252 100 6 Q
port 3 nsew signal output
rlabel metal2 s 243 93 253 99 6 Q
port 3 nsew signal output
rlabel metal1 s 243 16 248 140 6 Q
port 3 nsew signal output
rlabel metal1 s 243 92 252 100 6 Q
port 3 nsew signal output
rlabel metal1 s 243 93 253 100 6 Q
port 3 nsew signal output
rlabel metal2 s 229 79 237 87 6 QN
port 4 nsew signal output
rlabel metal2 s 228 80 238 86 6 QN
port 4 nsew signal output
rlabel metal1 s 209 16 214 43 6 QN
port 4 nsew signal output
rlabel metal1 s 209 80 214 140 6 QN
port 4 nsew signal output
rlabel metal1 s 209 38 236 43 6 QN
port 4 nsew signal output
rlabel metal1 s 231 38 236 86 6 QN
port 4 nsew signal output
rlabel metal1 s 209 80 238 86 6 QN
port 4 nsew signal output
rlabel metal2 s 10 147 18 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 34 147 42 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 33 148 43 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 58 147 66 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 57 148 67 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 82 147 90 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 81 148 91 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 106 147 114 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 105 148 115 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 130 147 138 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 129 148 139 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 154 147 162 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 153 148 163 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 178 147 186 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 177 148 187 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 202 147 210 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 201 148 211 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 226 147 234 155 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 225 148 235 154 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 28 106 33 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 89 106 94 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 145 121 150 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 177 106 182 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 226 106 231 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 0 147 260 159 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 34 1 42 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 33 2 43 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 58 1 66 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 57 2 67 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 82 1 90 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 81 2 91 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 106 1 114 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 105 2 115 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 130 1 138 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 129 2 139 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 154 1 162 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 153 2 163 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 178 1 186 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 177 2 187 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 202 1 210 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 201 2 211 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 226 1 234 9 6 VSS
port 6 nsew ground bidirectional
rlabel metal2 s 225 2 235 8 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 28 -3 33 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 89 -3 94 25 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 145 -3 150 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 177 -3 182 26 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 226 -3 231 33 6 VSS
port 6 nsew ground bidirectional
rlabel metal1 s 0 -3 260 9 6 VSS
port 6 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 -3 260 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
