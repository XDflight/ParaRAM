magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< ndiff >>
rect -42 399 42 418
rect -42 -399 -23 399
rect 23 -399 42 399
rect -42 -418 42 -399
<< ndiffc >>
rect -23 -399 23 399
<< metal1 >>
rect -34 399 34 410
rect -34 -399 -23 399
rect 23 -399 34 399
rect -34 -410 34 -399
<< properties >>
string GDS_END 325836
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 325064
<< end >>
