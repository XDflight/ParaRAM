magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 454 89 526
rect 193 454 313 526
rect 417 454 537 526
rect 641 454 761 526
rect -31 -73 89 -1
rect 193 -73 313 -1
rect 417 -73 537 -1
rect 641 -73 761 -1
use nmos_5p04310591302012_512x8m81  nmos_5p04310591302012_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 880 498
<< properties >>
string GDS_END 356816
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 356182
<< end >>
