magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 2344 938
<< mvpmos >>
rect 0 0 120 818
rect 224 0 344 818
rect 448 0 568 818
rect 672 0 792 818
rect 896 0 1016 818
rect 1120 0 1240 818
rect 1344 0 1464 818
rect 1568 0 1688 818
rect 1792 0 1912 818
rect 2016 0 2136 818
<< mvpdiff >>
rect -88 805 0 818
rect -88 759 -75 805
rect -29 759 0 805
rect -88 699 0 759
rect -88 653 -75 699
rect -29 653 0 699
rect -88 593 0 653
rect -88 547 -75 593
rect -29 547 0 593
rect -88 487 0 547
rect -88 441 -75 487
rect -29 441 0 487
rect -88 380 0 441
rect -88 334 -75 380
rect -29 334 0 380
rect -88 273 0 334
rect -88 227 -75 273
rect -29 227 0 273
rect -88 166 0 227
rect -88 120 -75 166
rect -29 120 0 166
rect -88 59 0 120
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 805 224 818
rect 120 759 149 805
rect 195 759 224 805
rect 120 699 224 759
rect 120 653 149 699
rect 195 653 224 699
rect 120 593 224 653
rect 120 547 149 593
rect 195 547 224 593
rect 120 487 224 547
rect 120 441 149 487
rect 195 441 224 487
rect 120 380 224 441
rect 120 334 149 380
rect 195 334 224 380
rect 120 273 224 334
rect 120 227 149 273
rect 195 227 224 273
rect 120 166 224 227
rect 120 120 149 166
rect 195 120 224 166
rect 120 59 224 120
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 805 448 818
rect 344 759 373 805
rect 419 759 448 805
rect 344 699 448 759
rect 344 653 373 699
rect 419 653 448 699
rect 344 593 448 653
rect 344 547 373 593
rect 419 547 448 593
rect 344 487 448 547
rect 344 441 373 487
rect 419 441 448 487
rect 344 380 448 441
rect 344 334 373 380
rect 419 334 448 380
rect 344 273 448 334
rect 344 227 373 273
rect 419 227 448 273
rect 344 166 448 227
rect 344 120 373 166
rect 419 120 448 166
rect 344 59 448 120
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 805 672 818
rect 568 759 597 805
rect 643 759 672 805
rect 568 699 672 759
rect 568 653 597 699
rect 643 653 672 699
rect 568 593 672 653
rect 568 547 597 593
rect 643 547 672 593
rect 568 487 672 547
rect 568 441 597 487
rect 643 441 672 487
rect 568 380 672 441
rect 568 334 597 380
rect 643 334 672 380
rect 568 273 672 334
rect 568 227 597 273
rect 643 227 672 273
rect 568 166 672 227
rect 568 120 597 166
rect 643 120 672 166
rect 568 59 672 120
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 805 896 818
rect 792 759 821 805
rect 867 759 896 805
rect 792 699 896 759
rect 792 653 821 699
rect 867 653 896 699
rect 792 593 896 653
rect 792 547 821 593
rect 867 547 896 593
rect 792 487 896 547
rect 792 441 821 487
rect 867 441 896 487
rect 792 380 896 441
rect 792 334 821 380
rect 867 334 896 380
rect 792 273 896 334
rect 792 227 821 273
rect 867 227 896 273
rect 792 166 896 227
rect 792 120 821 166
rect 867 120 896 166
rect 792 59 896 120
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 805 1120 818
rect 1016 759 1045 805
rect 1091 759 1120 805
rect 1016 699 1120 759
rect 1016 653 1045 699
rect 1091 653 1120 699
rect 1016 593 1120 653
rect 1016 547 1045 593
rect 1091 547 1120 593
rect 1016 487 1120 547
rect 1016 441 1045 487
rect 1091 441 1120 487
rect 1016 380 1120 441
rect 1016 334 1045 380
rect 1091 334 1120 380
rect 1016 273 1120 334
rect 1016 227 1045 273
rect 1091 227 1120 273
rect 1016 166 1120 227
rect 1016 120 1045 166
rect 1091 120 1120 166
rect 1016 59 1120 120
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 805 1344 818
rect 1240 759 1269 805
rect 1315 759 1344 805
rect 1240 699 1344 759
rect 1240 653 1269 699
rect 1315 653 1344 699
rect 1240 593 1344 653
rect 1240 547 1269 593
rect 1315 547 1344 593
rect 1240 487 1344 547
rect 1240 441 1269 487
rect 1315 441 1344 487
rect 1240 380 1344 441
rect 1240 334 1269 380
rect 1315 334 1344 380
rect 1240 273 1344 334
rect 1240 227 1269 273
rect 1315 227 1344 273
rect 1240 166 1344 227
rect 1240 120 1269 166
rect 1315 120 1344 166
rect 1240 59 1344 120
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 805 1568 818
rect 1464 759 1493 805
rect 1539 759 1568 805
rect 1464 699 1568 759
rect 1464 653 1493 699
rect 1539 653 1568 699
rect 1464 593 1568 653
rect 1464 547 1493 593
rect 1539 547 1568 593
rect 1464 487 1568 547
rect 1464 441 1493 487
rect 1539 441 1568 487
rect 1464 380 1568 441
rect 1464 334 1493 380
rect 1539 334 1568 380
rect 1464 273 1568 334
rect 1464 227 1493 273
rect 1539 227 1568 273
rect 1464 166 1568 227
rect 1464 120 1493 166
rect 1539 120 1568 166
rect 1464 59 1568 120
rect 1464 13 1493 59
rect 1539 13 1568 59
rect 1464 0 1568 13
rect 1688 805 1792 818
rect 1688 759 1717 805
rect 1763 759 1792 805
rect 1688 699 1792 759
rect 1688 653 1717 699
rect 1763 653 1792 699
rect 1688 593 1792 653
rect 1688 547 1717 593
rect 1763 547 1792 593
rect 1688 487 1792 547
rect 1688 441 1717 487
rect 1763 441 1792 487
rect 1688 380 1792 441
rect 1688 334 1717 380
rect 1763 334 1792 380
rect 1688 273 1792 334
rect 1688 227 1717 273
rect 1763 227 1792 273
rect 1688 166 1792 227
rect 1688 120 1717 166
rect 1763 120 1792 166
rect 1688 59 1792 120
rect 1688 13 1717 59
rect 1763 13 1792 59
rect 1688 0 1792 13
rect 1912 805 2016 818
rect 1912 759 1941 805
rect 1987 759 2016 805
rect 1912 699 2016 759
rect 1912 653 1941 699
rect 1987 653 2016 699
rect 1912 593 2016 653
rect 1912 547 1941 593
rect 1987 547 2016 593
rect 1912 487 2016 547
rect 1912 441 1941 487
rect 1987 441 2016 487
rect 1912 380 2016 441
rect 1912 334 1941 380
rect 1987 334 2016 380
rect 1912 273 2016 334
rect 1912 227 1941 273
rect 1987 227 2016 273
rect 1912 166 2016 227
rect 1912 120 1941 166
rect 1987 120 2016 166
rect 1912 59 2016 120
rect 1912 13 1941 59
rect 1987 13 2016 59
rect 1912 0 2016 13
rect 2136 805 2224 818
rect 2136 759 2165 805
rect 2211 759 2224 805
rect 2136 699 2224 759
rect 2136 653 2165 699
rect 2211 653 2224 699
rect 2136 593 2224 653
rect 2136 547 2165 593
rect 2211 547 2224 593
rect 2136 487 2224 547
rect 2136 441 2165 487
rect 2211 441 2224 487
rect 2136 380 2224 441
rect 2136 334 2165 380
rect 2211 334 2224 380
rect 2136 273 2224 334
rect 2136 227 2165 273
rect 2211 227 2224 273
rect 2136 166 2224 227
rect 2136 120 2165 166
rect 2211 120 2224 166
rect 2136 59 2224 120
rect 2136 13 2165 59
rect 2211 13 2224 59
rect 2136 0 2224 13
<< mvpdiffc >>
rect -75 759 -29 805
rect -75 653 -29 699
rect -75 547 -29 593
rect -75 441 -29 487
rect -75 334 -29 380
rect -75 227 -29 273
rect -75 120 -29 166
rect -75 13 -29 59
rect 149 759 195 805
rect 149 653 195 699
rect 149 547 195 593
rect 149 441 195 487
rect 149 334 195 380
rect 149 227 195 273
rect 149 120 195 166
rect 149 13 195 59
rect 373 759 419 805
rect 373 653 419 699
rect 373 547 419 593
rect 373 441 419 487
rect 373 334 419 380
rect 373 227 419 273
rect 373 120 419 166
rect 373 13 419 59
rect 597 759 643 805
rect 597 653 643 699
rect 597 547 643 593
rect 597 441 643 487
rect 597 334 643 380
rect 597 227 643 273
rect 597 120 643 166
rect 597 13 643 59
rect 821 759 867 805
rect 821 653 867 699
rect 821 547 867 593
rect 821 441 867 487
rect 821 334 867 380
rect 821 227 867 273
rect 821 120 867 166
rect 821 13 867 59
rect 1045 759 1091 805
rect 1045 653 1091 699
rect 1045 547 1091 593
rect 1045 441 1091 487
rect 1045 334 1091 380
rect 1045 227 1091 273
rect 1045 120 1091 166
rect 1045 13 1091 59
rect 1269 759 1315 805
rect 1269 653 1315 699
rect 1269 547 1315 593
rect 1269 441 1315 487
rect 1269 334 1315 380
rect 1269 227 1315 273
rect 1269 120 1315 166
rect 1269 13 1315 59
rect 1493 759 1539 805
rect 1493 653 1539 699
rect 1493 547 1539 593
rect 1493 441 1539 487
rect 1493 334 1539 380
rect 1493 227 1539 273
rect 1493 120 1539 166
rect 1493 13 1539 59
rect 1717 759 1763 805
rect 1717 653 1763 699
rect 1717 547 1763 593
rect 1717 441 1763 487
rect 1717 334 1763 380
rect 1717 227 1763 273
rect 1717 120 1763 166
rect 1717 13 1763 59
rect 1941 759 1987 805
rect 1941 653 1987 699
rect 1941 547 1987 593
rect 1941 441 1987 487
rect 1941 334 1987 380
rect 1941 227 1987 273
rect 1941 120 1987 166
rect 1941 13 1987 59
rect 2165 759 2211 805
rect 2165 653 2211 699
rect 2165 547 2211 593
rect 2165 441 2211 487
rect 2165 334 2211 380
rect 2165 227 2211 273
rect 2165 120 2211 166
rect 2165 13 2211 59
<< polysilicon >>
rect 0 818 120 862
rect 224 818 344 862
rect 448 818 568 862
rect 672 818 792 862
rect 896 818 1016 862
rect 1120 818 1240 862
rect 1344 818 1464 862
rect 1568 818 1688 862
rect 1792 818 1912 862
rect 2016 818 2136 862
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
<< metal1 >>
rect -75 805 -29 818
rect -75 699 -29 759
rect -75 593 -29 653
rect -75 487 -29 547
rect -75 380 -29 441
rect -75 273 -29 334
rect -75 166 -29 227
rect -75 59 -29 120
rect -75 0 -29 13
rect 149 805 195 818
rect 149 699 195 759
rect 149 593 195 653
rect 149 487 195 547
rect 149 380 195 441
rect 149 273 195 334
rect 149 166 195 227
rect 149 59 195 120
rect 149 0 195 13
rect 373 805 419 818
rect 373 699 419 759
rect 373 593 419 653
rect 373 487 419 547
rect 373 380 419 441
rect 373 273 419 334
rect 373 166 419 227
rect 373 59 419 120
rect 373 0 419 13
rect 597 805 643 818
rect 597 699 643 759
rect 597 593 643 653
rect 597 487 643 547
rect 597 380 643 441
rect 597 273 643 334
rect 597 166 643 227
rect 597 59 643 120
rect 597 0 643 13
rect 821 805 867 818
rect 821 699 867 759
rect 821 593 867 653
rect 821 487 867 547
rect 821 380 867 441
rect 821 273 867 334
rect 821 166 867 227
rect 821 59 867 120
rect 821 0 867 13
rect 1045 805 1091 818
rect 1045 699 1091 759
rect 1045 593 1091 653
rect 1045 487 1091 547
rect 1045 380 1091 441
rect 1045 273 1091 334
rect 1045 166 1091 227
rect 1045 59 1091 120
rect 1045 0 1091 13
rect 1269 805 1315 818
rect 1269 699 1315 759
rect 1269 593 1315 653
rect 1269 487 1315 547
rect 1269 380 1315 441
rect 1269 273 1315 334
rect 1269 166 1315 227
rect 1269 59 1315 120
rect 1269 0 1315 13
rect 1493 805 1539 818
rect 1493 699 1539 759
rect 1493 593 1539 653
rect 1493 487 1539 547
rect 1493 380 1539 441
rect 1493 273 1539 334
rect 1493 166 1539 227
rect 1493 59 1539 120
rect 1493 0 1539 13
rect 1717 805 1763 818
rect 1717 699 1763 759
rect 1717 593 1763 653
rect 1717 487 1763 547
rect 1717 380 1763 441
rect 1717 273 1763 334
rect 1717 166 1763 227
rect 1717 59 1763 120
rect 1717 0 1763 13
rect 1941 805 1987 818
rect 1941 699 1987 759
rect 1941 593 1987 653
rect 1941 487 1987 547
rect 1941 380 1987 441
rect 1941 273 1987 334
rect 1941 166 1987 227
rect 1941 59 1987 120
rect 1941 0 1987 13
rect 2165 805 2211 818
rect 2165 699 2211 759
rect 2165 593 2211 653
rect 2165 487 2211 547
rect 2165 380 2211 441
rect 2165 273 2211 334
rect 2165 166 2211 227
rect 2165 59 2211 120
rect 2165 0 2211 13
<< labels >>
flabel metal1 s -52 409 -52 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 2188 409 2188 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 409 172 409 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 409 396 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 409 620 409 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 409 844 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 409 1068 409 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 409 1292 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 409 1516 409 0 FreeSans 400 0 0 0 D
flabel metal1 s 1740 409 1740 409 0 FreeSans 400 0 0 0 S
flabel metal1 s 1964 409 1964 409 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 56090
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 46060
<< end >>
