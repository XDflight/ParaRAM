magic
tech gf180mcuB
timestamp 1666464484
<< metal1 >>
rect 0 111 82 123
rect 11 70 16 111
rect 45 70 54 111
rect 66 77 71 104
rect 66 76 74 77
rect 66 70 76 76
rect 66 69 74 70
rect 39 57 49 63
rect 12 44 22 50
rect 42 12 54 36
rect 66 19 71 69
rect 0 0 82 12
<< obsm1 >>
rect 28 50 33 104
rect 55 50 61 52
rect 28 44 61 50
rect 28 34 33 44
rect 55 42 61 44
rect 14 29 33 34
rect 14 19 19 29
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 66 69 76 77
rect 39 56 49 64
rect 13 50 21 51
rect 12 44 22 50
rect 13 43 21 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 s 13 43 21 51 6 A
port 1 nsew signal input
rlabel metal2 s 12 44 22 50 6 A
port 1 nsew signal input
rlabel metal1 s 12 44 22 50 6 A
port 1 nsew signal input
rlabel metal2 s 39 56 49 64 6 B
port 2 nsew signal input
rlabel metal1 s 39 57 49 63 6 B
port 2 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 45 70 54 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 111 82 123 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 42 0 54 36 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 0 0 82 12 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 66 69 76 77 6 Y
port 5 nsew signal output
rlabel metal1 s 66 19 71 104 6 Y
port 5 nsew signal output
rlabel metal1 s 66 69 74 77 6 Y
port 5 nsew signal output
rlabel metal1 s 66 70 76 76 6 Y
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 82 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
