magic
tech gf180mcuB
magscale 1 5
timestamp 1667403392
<< checkpaint >>
rect 15600 15600 36500 36500
<< metal4 >>
rect 16600 27040 18100 35500
tri 18100 27040 18722 27662 sw
tri 16600 25088 18552 27040 ne
rect 18552 25088 18722 27040
tri 18722 25088 20674 27040 sw
tri 18552 22966 20674 25088 ne
tri 20674 22966 22796 25088 sw
tri 20674 20844 22796 22966 ne
tri 22796 20844 24918 22966 sw
tri 22796 18722 24918 20844 ne
tri 24918 18722 27040 20844 sw
tri 24918 16600 27040 18722 ne
tri 27040 18100 27662 18722 sw
rect 27040 16600 35500 18100
<< end >>
