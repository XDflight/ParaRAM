magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 344 1275
<< polysilicon >>
rect -31 1134 89 1206
rect -31 -74 89 -1
use pmos_5p04310589983264_64x8m81  pmos_5p04310589983264_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 1254
<< properties >>
string GDS_END 140908
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 140594
<< end >>
