magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -3742 323 3742 342
rect -3742 -323 -3723 323
rect 3723 -323 3742 323
rect -3742 -342 3742 -323
<< psubdiffcont >>
rect -3723 -323 3723 323
<< metal1 >>
rect -3734 323 3734 334
rect -3734 -323 -3723 323
rect 3723 -323 3734 323
rect -3734 -334 3734 -323
<< properties >>
string GDS_END 701796
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 668000
<< end >>
