magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 822
<< mvpmos >>
rect 0 0 120 702
rect 224 0 344 702
<< mvpdiff >>
rect -88 689 0 702
rect -88 643 -75 689
rect -29 643 0 689
rect -88 584 0 643
rect -88 538 -75 584
rect -29 538 0 584
rect -88 479 0 538
rect -88 433 -75 479
rect -29 433 0 479
rect -88 374 0 433
rect -88 328 -75 374
rect -29 328 0 374
rect -88 269 0 328
rect -88 223 -75 269
rect -29 223 0 269
rect -88 164 0 223
rect -88 118 -75 164
rect -29 118 0 164
rect -88 59 0 118
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 689 224 702
rect 120 643 149 689
rect 195 643 224 689
rect 120 584 224 643
rect 120 538 149 584
rect 195 538 224 584
rect 120 479 224 538
rect 120 433 149 479
rect 195 433 224 479
rect 120 374 224 433
rect 120 328 149 374
rect 195 328 224 374
rect 120 269 224 328
rect 120 223 149 269
rect 195 223 224 269
rect 120 164 224 223
rect 120 118 149 164
rect 195 118 224 164
rect 120 59 224 118
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 689 432 702
rect 344 643 373 689
rect 419 643 432 689
rect 344 584 432 643
rect 344 538 373 584
rect 419 538 432 584
rect 344 479 432 538
rect 344 433 373 479
rect 419 433 432 479
rect 344 374 432 433
rect 344 328 373 374
rect 419 328 432 374
rect 344 269 432 328
rect 344 223 373 269
rect 419 223 432 269
rect 344 164 432 223
rect 344 118 373 164
rect 419 118 432 164
rect 344 59 432 118
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 643 -29 689
rect -75 538 -29 584
rect -75 433 -29 479
rect -75 328 -29 374
rect -75 223 -29 269
rect -75 118 -29 164
rect -75 13 -29 59
rect 149 643 195 689
rect 149 538 195 584
rect 149 433 195 479
rect 149 328 195 374
rect 149 223 195 269
rect 149 118 195 164
rect 149 13 195 59
rect 373 643 419 689
rect 373 538 419 584
rect 373 433 419 479
rect 373 328 419 374
rect 373 223 419 269
rect 373 118 419 164
rect 373 13 419 59
<< polysilicon >>
rect 0 702 120 746
rect 224 702 344 746
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 689 -29 702
rect -75 584 -29 643
rect -75 479 -29 538
rect -75 374 -29 433
rect -75 269 -29 328
rect -75 164 -29 223
rect -75 59 -29 118
rect -75 0 -29 13
rect 149 689 195 702
rect 149 584 195 643
rect 149 479 195 538
rect 149 374 195 433
rect 149 269 195 328
rect 149 164 195 223
rect 149 59 195 118
rect 149 0 195 13
rect 373 689 419 702
rect 373 584 419 643
rect 373 479 419 538
rect 373 374 419 433
rect 373 269 419 328
rect 373 164 419 223
rect 373 59 419 118
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 351 -52 351 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 351 396 351 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 351 172 351 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 1108358
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1105672
<< end >>
