magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 3446 1094
<< pwell >>
rect -86 -86 3446 453
<< mvnmos >>
rect 124 175 244 333
rect 348 175 468 333
rect 716 156 836 274
rect 940 156 1060 274
rect 1164 156 1284 274
rect 1332 156 1452 274
rect 1644 215 1764 333
rect 1868 215 1988 333
rect 2092 215 2212 333
rect 2360 175 2480 333
rect 2672 175 2792 333
rect 3040 69 3160 333
<< mvpmos >>
rect 144 573 244 849
rect 348 573 448 849
rect 736 592 836 792
rect 960 592 1060 792
rect 1164 592 1264 792
rect 1352 592 1452 792
rect 1644 592 1744 792
rect 1868 592 1968 792
rect 2120 592 2220 792
rect 2380 631 2480 851
rect 2612 631 2712 851
rect 3040 573 3140 939
<< mvndiff >>
rect 36 320 124 333
rect 36 274 49 320
rect 95 274 124 320
rect 36 175 124 274
rect 244 234 348 333
rect 244 188 273 234
rect 319 188 348 234
rect 244 175 348 188
rect 468 320 556 333
rect 468 274 497 320
rect 543 274 556 320
rect 1564 274 1644 333
rect 468 175 556 274
rect 628 215 716 274
rect 628 169 641 215
rect 687 169 716 215
rect 628 156 716 169
rect 836 261 940 274
rect 836 215 865 261
rect 911 215 940 261
rect 836 156 940 215
rect 1060 261 1164 274
rect 1060 215 1089 261
rect 1135 215 1164 261
rect 1060 156 1164 215
rect 1284 156 1332 274
rect 1452 215 1644 274
rect 1764 320 1868 333
rect 1764 274 1793 320
rect 1839 274 1868 320
rect 1764 215 1868 274
rect 1988 320 2092 333
rect 1988 274 2017 320
rect 2063 274 2092 320
rect 1988 215 2092 274
rect 2212 234 2360 333
rect 2212 215 2285 234
rect 1452 156 1584 215
rect 1512 114 1584 156
rect 2272 188 2285 215
rect 2331 188 2360 234
rect 2272 175 2360 188
rect 2480 175 2672 333
rect 2792 320 2880 333
rect 2792 274 2821 320
rect 2867 274 2880 320
rect 2792 175 2880 274
rect 2952 320 3040 333
rect 2952 274 2965 320
rect 3011 274 3040 320
rect 1512 68 1525 114
rect 1571 68 1584 114
rect 1512 55 1584 68
rect 2540 114 2612 175
rect 2540 68 2553 114
rect 2599 68 2612 114
rect 2952 69 3040 274
rect 3160 222 3248 333
rect 3160 82 3189 222
rect 3235 82 3248 222
rect 3160 69 3248 82
rect 2540 55 2612 68
<< mvpdiff >>
rect 56 739 144 849
rect 56 599 69 739
rect 115 599 144 739
rect 56 573 144 599
rect 244 836 348 849
rect 244 696 273 836
rect 319 696 348 836
rect 244 573 348 696
rect 448 632 536 849
rect 2300 792 2380 851
rect 448 586 477 632
rect 523 586 536 632
rect 648 779 736 792
rect 648 733 661 779
rect 707 733 736 779
rect 648 592 736 733
rect 836 745 960 792
rect 836 605 885 745
rect 931 605 960 745
rect 836 592 960 605
rect 1060 745 1164 792
rect 1060 605 1089 745
rect 1135 605 1164 745
rect 1060 592 1164 605
rect 1264 592 1352 792
rect 1452 779 1644 792
rect 1452 639 1481 779
rect 1527 639 1644 779
rect 1452 592 1644 639
rect 1744 745 1868 792
rect 1744 605 1793 745
rect 1839 605 1868 745
rect 1744 592 1868 605
rect 1968 745 2120 792
rect 1968 605 2017 745
rect 2063 605 2120 745
rect 1968 592 2120 605
rect 2220 735 2380 792
rect 2220 689 2305 735
rect 2351 689 2380 735
rect 2220 631 2380 689
rect 2480 838 2612 851
rect 2480 792 2509 838
rect 2555 792 2612 838
rect 2480 631 2612 792
rect 2712 632 2844 851
rect 2712 631 2785 632
rect 2220 592 2300 631
rect 448 573 536 586
rect 2772 586 2785 631
rect 2831 586 2844 632
rect 2772 573 2844 586
rect 2952 632 3040 939
rect 2952 586 2965 632
rect 3011 586 3040 632
rect 2952 573 3040 586
rect 3140 926 3228 939
rect 3140 786 3169 926
rect 3215 786 3228 926
rect 3140 573 3228 786
<< mvndiffc >>
rect 49 274 95 320
rect 273 188 319 234
rect 497 274 543 320
rect 641 169 687 215
rect 865 215 911 261
rect 1089 215 1135 261
rect 1793 274 1839 320
rect 2017 274 2063 320
rect 2285 188 2331 234
rect 2821 274 2867 320
rect 2965 274 3011 320
rect 1525 68 1571 114
rect 2553 68 2599 114
rect 3189 82 3235 222
<< mvpdiffc >>
rect 69 599 115 739
rect 273 696 319 836
rect 477 586 523 632
rect 661 733 707 779
rect 885 605 931 745
rect 1089 605 1135 745
rect 1481 639 1527 779
rect 1793 605 1839 745
rect 2017 605 2063 745
rect 2305 689 2351 735
rect 2509 792 2555 838
rect 2785 586 2831 632
rect 2965 586 3011 632
rect 3169 786 3215 926
<< polysilicon >>
rect 348 909 1060 949
rect 3040 939 3140 983
rect 144 849 244 893
rect 348 849 448 909
rect 736 792 836 836
rect 960 792 1060 909
rect 1164 884 1968 924
rect 1164 871 1264 884
rect 1164 825 1177 871
rect 1223 825 1264 871
rect 1164 792 1264 825
rect 1352 792 1452 836
rect 1644 792 1744 836
rect 1868 792 1968 884
rect 2380 851 2480 895
rect 2612 851 2712 895
rect 2120 792 2220 836
rect 144 504 244 573
rect 144 458 157 504
rect 203 458 244 504
rect 144 377 244 458
rect 124 333 244 377
rect 348 412 448 573
rect 348 366 361 412
rect 407 377 448 412
rect 736 512 836 592
rect 960 548 1060 592
rect 736 466 777 512
rect 823 466 836 512
rect 1164 500 1264 592
rect 407 366 468 377
rect 348 333 468 366
rect 736 318 836 466
rect 1020 460 1264 500
rect 1352 559 1452 592
rect 1352 513 1393 559
rect 1439 513 1452 559
rect 1020 318 1060 460
rect 716 274 836 318
rect 940 274 1060 318
rect 1164 353 1284 366
rect 1164 307 1225 353
rect 1271 307 1284 353
rect 1352 318 1452 513
rect 1644 445 1744 592
rect 1868 500 1968 592
rect 2120 548 2220 592
rect 2180 519 2220 548
rect 2180 506 2252 519
rect 1868 460 2132 500
rect 1644 399 1657 445
rect 1703 399 1744 445
rect 1644 377 1744 399
rect 2092 377 2132 460
rect 2180 460 2193 506
rect 2239 460 2252 506
rect 2180 447 2252 460
rect 2380 492 2480 631
rect 2380 446 2421 492
rect 2467 446 2480 492
rect 2380 377 2480 446
rect 2612 598 2712 631
rect 2612 552 2625 598
rect 2671 552 2712 598
rect 2612 393 2712 552
rect 3040 482 3140 573
rect 2837 469 3140 482
rect 2837 423 2850 469
rect 2896 423 3140 469
rect 2837 410 3140 423
rect 1644 333 1764 377
rect 1868 333 1988 377
rect 2092 333 2212 377
rect 2360 333 2480 377
rect 2672 333 2792 393
rect 3040 377 3140 410
rect 3040 333 3160 377
rect 1164 274 1284 307
rect 1332 274 1452 318
rect 124 131 244 175
rect 348 64 468 175
rect 1644 171 1764 215
rect 1868 182 1988 215
rect 716 112 836 156
rect 940 112 1060 156
rect 1164 64 1284 156
rect 1332 112 1452 156
rect 1868 136 1881 182
rect 1927 136 1988 182
rect 2092 171 2212 215
rect 1868 123 1988 136
rect 2360 131 2480 175
rect 348 24 1284 64
rect 2672 131 2792 175
rect 3040 25 3160 69
<< polycontact >>
rect 1177 825 1223 871
rect 157 458 203 504
rect 361 366 407 412
rect 777 466 823 512
rect 1393 513 1439 559
rect 1225 307 1271 353
rect 1657 399 1703 445
rect 2193 460 2239 506
rect 2421 446 2467 492
rect 2625 552 2671 598
rect 2850 423 2896 469
rect 1881 136 1927 182
<< metal1 >>
rect 0 926 3360 1098
rect 0 918 3169 926
rect 273 836 319 918
rect 69 739 115 750
rect 661 779 707 918
rect 661 722 707 733
rect 753 825 1177 871
rect 1223 825 1234 871
rect 273 685 319 696
rect 753 644 799 825
rect 1481 779 1527 918
rect 2509 838 2555 918
rect 2509 781 2555 792
rect 3215 918 3360 926
rect 115 599 407 634
rect 69 588 407 599
rect 142 504 314 542
rect 142 458 157 504
rect 203 458 314 504
rect 142 447 314 458
rect 361 412 407 588
rect 361 348 407 366
rect 49 320 407 348
rect 95 302 407 320
rect 477 632 799 644
rect 523 598 799 632
rect 885 745 958 756
rect 931 605 958 745
rect 523 586 543 598
rect 885 594 958 605
rect 477 320 543 586
rect 690 512 866 542
rect 690 466 777 512
rect 823 466 866 512
rect 49 263 95 274
rect 477 274 497 320
rect 477 263 543 274
rect 912 272 958 594
rect 865 261 958 272
rect 273 234 319 245
rect 273 90 319 188
rect 641 215 687 226
rect 911 215 958 261
rect 865 204 958 215
rect 1089 745 1135 756
rect 3169 775 3215 786
rect 1481 628 1527 639
rect 1793 745 1839 756
rect 1089 456 1135 605
rect 1793 570 1839 605
rect 1393 559 1839 570
rect 1439 513 1839 559
rect 1393 502 1839 513
rect 1089 445 1703 456
rect 1089 410 1657 445
rect 1089 261 1135 410
rect 1657 388 1703 399
rect 1089 204 1135 215
rect 1225 353 1271 364
rect 1225 217 1271 307
rect 1793 320 1839 502
rect 1793 263 1839 274
rect 2017 745 2063 756
rect 2294 689 2305 735
rect 2351 689 3103 735
rect 2017 598 2063 605
rect 2785 632 2831 643
rect 2017 552 2625 598
rect 2671 552 2682 598
rect 2017 320 2063 552
rect 2017 263 2063 274
rect 2109 460 2193 506
rect 2239 460 2250 506
rect 2785 492 2831 586
rect 2109 217 2155 460
rect 2410 446 2421 492
rect 2467 491 2831 492
rect 2942 632 3011 643
rect 2942 586 2965 632
rect 2467 469 2896 491
rect 2467 446 2850 469
rect 2821 423 2850 446
rect 2821 320 2896 423
rect 2867 274 2896 320
rect 2821 263 2896 274
rect 2942 320 3011 586
rect 2942 274 2965 320
rect 2942 263 3011 274
rect 1225 182 2155 217
rect 1225 171 1881 182
rect 641 90 687 169
rect 1870 136 1881 171
rect 1927 136 2155 182
rect 2285 234 2331 245
rect 3057 217 3103 689
rect 2331 188 3103 217
rect 2285 171 3103 188
rect 3189 222 3235 233
rect 1525 114 1571 125
rect 0 68 1525 90
rect 2553 114 2599 125
rect 1571 68 2553 90
rect 2599 82 3189 90
rect 3235 82 3360 90
rect 2599 68 3360 82
rect 0 -90 3360 68
<< labels >>
flabel metal1 s 142 447 314 542 0 FreeSans 200 0 0 0 CLKN
port 2 nsew clock input
flabel metal1 s 690 466 866 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 2942 263 3011 643 0 FreeSans 200 0 0 0 Q
port 3 nsew default output
flabel metal1 s 0 918 3360 1098 0 FreeSans 200 0 0 0 VDD
port 4 nsew power bidirectional abutment
flabel metal1 s 273 233 319 245 0 FreeSans 200 0 0 0 VSS
port 7 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3169 781 3215 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 2509 781 2555 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1481 781 1527 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 661 781 707 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 781 319 918 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3169 775 3215 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1481 775 1527 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 661 775 707 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 781 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1481 722 1527 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 661 722 707 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 722 319 775 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1481 685 1527 722 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 273 685 319 722 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1481 628 1527 685 1 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 3189 226 3235 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 226 319 233 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3189 125 3235 226 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 641 125 687 226 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 226 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 3189 90 3235 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 2553 90 2599 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1525 90 1571 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 641 90 687 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 125 1 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3360 90 1 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 1008
string GDS_END 1464828
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1457334
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
