magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect 0 459 112 549
rect 0 -45 112 45
<< labels >>
rlabel metal1 s 0 459 112 549 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -45 112 45 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 112 504
string GDS_END 753040
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 752006
string LEFclass core SPACER
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
