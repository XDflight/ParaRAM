magic
tech gf180mcuA
timestamp 1667403424
<< metal1 >>
rect -81 147 293 159
rect -70 106 -65 147
rect -70 93 -60 99
rect -4 121 1 147
rect 28 106 33 147
rect 89 106 94 147
rect 145 121 150 147
rect -13 80 -3 86
rect 52 80 75 86
rect 38 67 48 73
rect 67 47 73 80
rect 194 131 199 147
rect 110 80 131 86
rect -70 9 -65 33
rect -35 9 -30 33
rect 65 41 75 47
rect 110 46 116 80
rect 153 80 163 86
rect 198 80 208 86
rect 243 86 248 140
rect 260 106 265 147
rect 277 100 282 140
rect 277 93 287 100
rect 277 92 286 93
rect 243 80 272 86
rect 108 40 118 46
rect 10 9 15 33
rect 28 9 33 33
rect 89 9 94 25
rect 145 9 150 33
rect 180 9 185 33
rect 265 43 270 80
rect 243 38 270 43
rect 225 9 230 33
rect 243 16 248 38
rect 260 9 265 33
rect 277 16 282 92
rect -81 -3 293 9
<< obsm1 >>
rect -53 47 -48 140
rect -38 52 -33 140
rect -21 116 -16 140
rect 13 116 18 140
rect -21 111 18 116
rect 61 101 66 140
rect 117 121 122 140
rect 99 116 122 121
rect 28 96 66 101
rect 28 73 33 96
rect 81 93 91 99
rect -28 67 -18 73
rect 7 67 33 73
rect -38 47 -13 52
rect 9 47 14 48
rect 28 47 33 67
rect 83 47 89 93
rect 99 71 104 116
rect 134 93 144 99
rect 162 97 167 140
rect 177 126 182 140
rect 211 126 216 140
rect 177 121 216 126
rect 180 99 186 101
rect 228 99 233 140
rect 98 66 104 71
rect -55 41 -45 47
rect -18 41 17 47
rect 28 42 48 47
rect -53 40 -47 41
rect -53 16 -48 40
rect -18 16 -13 41
rect 9 40 14 41
rect 40 33 48 42
rect 81 41 91 47
rect 98 34 103 66
rect 136 73 142 93
rect 162 92 173 97
rect 168 73 173 92
rect 180 93 236 99
rect 180 91 186 93
rect 135 67 145 73
rect 162 68 173 73
rect 121 54 131 60
rect 162 52 168 68
rect 228 60 233 93
rect 208 54 257 60
rect 40 28 66 33
rect 98 29 125 34
rect 61 16 66 28
rect 117 28 125 29
rect 117 16 122 28
rect 162 16 167 52
rect 178 40 188 46
rect 208 16 213 54
rect 218 40 228 46
<< metal2 >>
rect -71 154 -63 155
rect -47 154 -39 155
rect -23 154 -15 155
rect 1 154 9 155
rect 25 154 33 155
rect 49 154 57 155
rect 73 154 81 155
rect 97 154 105 155
rect 121 154 129 155
rect 145 154 153 155
rect 169 154 177 155
rect 193 154 201 155
rect 217 154 225 155
rect 241 154 249 155
rect 265 154 273 155
rect -72 148 -62 154
rect -48 148 -38 154
rect -24 148 -14 154
rect 0 148 10 154
rect 24 148 34 154
rect 48 148 58 154
rect 72 148 82 154
rect 96 148 106 154
rect 120 148 130 154
rect 144 148 154 154
rect 168 148 178 154
rect 192 148 202 154
rect 216 148 226 154
rect 240 148 250 154
rect 264 148 274 154
rect -71 147 -63 148
rect -47 147 -39 148
rect -23 147 -15 148
rect 1 147 9 148
rect 25 147 33 148
rect 49 147 57 148
rect 73 147 81 148
rect 97 147 105 148
rect 121 147 129 148
rect 145 147 153 148
rect 169 147 177 148
rect 193 147 201 148
rect 217 147 225 148
rect 241 147 249 148
rect 265 147 273 148
rect -11 106 206 112
rect -70 92 -60 100
rect -11 87 -5 106
rect 200 87 206 106
rect 278 99 286 100
rect 277 93 287 99
rect 278 92 286 93
rect -13 79 -3 87
rect 65 86 74 87
rect 121 86 131 87
rect 154 86 162 87
rect 65 80 163 86
rect 65 79 74 80
rect 121 79 131 80
rect 154 79 162 80
rect 198 79 208 87
rect 263 86 271 87
rect 262 80 272 86
rect 263 79 271 80
rect 38 66 48 74
rect -71 8 -63 9
rect -47 8 -39 9
rect -23 8 -15 9
rect 1 8 9 9
rect 25 8 33 9
rect 49 8 57 9
rect 73 8 81 9
rect 97 8 105 9
rect 121 8 129 9
rect 145 8 153 9
rect 169 8 177 9
rect 193 8 201 9
rect 217 8 225 9
rect 241 8 249 9
rect 265 8 273 9
rect -72 2 -62 8
rect -48 2 -38 8
rect -24 2 -14 8
rect 0 2 10 8
rect 24 2 34 8
rect 48 2 58 8
rect 72 2 82 8
rect 96 2 106 8
rect 120 2 130 8
rect 144 2 154 8
rect 168 2 178 8
rect 192 2 202 8
rect 216 2 226 8
rect 240 2 250 8
rect 264 2 274 8
rect -71 1 -63 2
rect -47 1 -39 2
rect -23 1 -15 2
rect 1 1 9 2
rect 25 1 33 2
rect 49 1 57 2
rect 73 1 81 2
rect 97 1 105 2
rect 121 1 129 2
rect 145 1 153 2
rect 169 1 177 2
rect 193 1 201 2
rect 217 1 225 2
rect 241 1 249 2
rect 265 1 273 2
<< obsm2 >>
rect 135 99 143 100
rect 179 99 187 100
rect 134 93 188 99
rect 135 92 143 93
rect 179 92 187 93
rect 226 92 236 100
rect -28 66 -18 74
rect 7 66 17 74
rect 136 73 144 74
rect 135 67 145 73
rect 136 66 144 67
rect -55 47 -45 48
rect -26 47 -20 66
rect 122 60 130 61
rect 161 60 169 61
rect 248 60 256 61
rect 121 54 171 60
rect 241 54 257 60
rect 122 53 130 54
rect 161 53 169 54
rect 248 53 256 54
rect -55 41 -20 47
rect -55 40 -45 41
rect -26 21 -20 41
rect 7 47 17 48
rect 82 47 90 48
rect 7 41 91 47
rect 7 40 17 41
rect 82 40 90 41
rect 178 39 188 47
rect 216 39 228 47
rect 116 34 124 35
rect 178 34 186 39
rect 115 28 186 34
rect 116 27 124 28
rect 216 21 222 39
rect -26 15 222 21
<< labels >>
rlabel metal2 s 65 79 74 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 121 79 131 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 154 79 162 87 6 CLK
port 1 nsew clock input
rlabel metal2 s 65 80 163 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 67 41 73 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 65 41 75 47 6 CLK
port 1 nsew clock input
rlabel metal1 s 52 80 75 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 110 40 116 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 108 40 118 46 6 CLK
port 1 nsew clock input
rlabel metal1 s 110 80 131 86 6 CLK
port 1 nsew clock input
rlabel metal1 s 153 80 163 86 6 CLK
port 1 nsew clock input
rlabel metal2 s 38 66 48 74 6 D
port 2 nsew signal input
rlabel metal1 s 38 67 48 73 6 D
port 2 nsew signal input
rlabel metal2 s 278 92 286 100 6 Q
port 3 nsew signal output
rlabel metal2 s 277 93 287 99 6 Q
port 3 nsew signal output
rlabel metal1 s 277 16 282 140 6 Q
port 3 nsew signal output
rlabel metal1 s 277 92 286 100 6 Q
port 3 nsew signal output
rlabel metal1 s 277 93 287 100 6 Q
port 3 nsew signal output
rlabel metal2 s 263 79 271 87 6 QN
port 4 nsew signal output
rlabel metal2 s 262 80 272 86 6 QN
port 4 nsew signal output
rlabel metal1 s 243 16 248 43 6 QN
port 4 nsew signal output
rlabel metal1 s 243 80 248 140 6 QN
port 4 nsew signal output
rlabel metal1 s 243 38 270 43 6 QN
port 4 nsew signal output
rlabel metal1 s 265 38 270 86 6 QN
port 4 nsew signal output
rlabel metal1 s 243 80 272 86 6 QN
port 4 nsew signal output
rlabel metal2 s -70 92 -60 100 4 RN
port 5 nsew signal input
rlabel metal1 s -70 93 -60 99 4 RN
port 5 nsew signal input
rlabel metal2 s -11 79 -5 112 4 SN
port 6 nsew signal output
rlabel metal2 s -13 79 -3 87 4 SN
port 6 nsew signal output
rlabel metal2 s 200 79 206 112 6 SN
port 6 nsew signal output
rlabel metal2 s -11 106 206 112 6 SN
port 6 nsew signal output
rlabel metal2 s 198 79 208 87 6 SN
port 6 nsew signal output
rlabel metal1 s -13 80 -3 86 4 SN
port 6 nsew signal output
rlabel metal1 s 198 80 208 86 6 SN
port 6 nsew signal output
rlabel metal2 s -71 147 -63 155 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -72 148 -62 154 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -47 147 -39 155 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -48 148 -38 154 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -23 147 -15 155 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -24 148 -14 154 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 1 147 9 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 0 148 10 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 25 147 33 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 24 148 34 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 49 147 57 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 48 148 58 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 73 147 81 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 72 148 82 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 97 147 105 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 96 148 106 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 121 147 129 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 120 148 130 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 145 147 153 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 144 148 154 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 169 147 177 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 168 148 178 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 193 147 201 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 192 148 202 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 217 147 225 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 216 148 226 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 241 147 249 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 240 148 250 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 265 147 273 155 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s 264 148 274 154 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s -70 106 -65 159 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s -4 121 1 159 4 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 28 106 33 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 89 106 94 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 145 121 150 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 194 131 199 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 260 106 265 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s -81 147 293 159 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal2 s -71 1 -63 9 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s -72 2 -62 8 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s -47 1 -39 9 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s -48 2 -38 8 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s -23 1 -15 9 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s -24 2 -14 8 4 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 1 1 9 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 0 2 10 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 25 1 33 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 24 2 34 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 49 1 57 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 48 2 58 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 73 1 81 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 72 2 82 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 97 1 105 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 96 2 106 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 121 1 129 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 120 2 130 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 145 1 153 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 144 2 154 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 169 1 177 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 168 2 178 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 193 1 201 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 192 2 202 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 217 1 225 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 216 2 226 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 241 1 249 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 240 2 250 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 265 1 273 9 6 VSS
port 8 nsew ground bidirectional
rlabel metal2 s 264 2 274 8 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s -70 -3 -65 33 4 VSS
port 8 nsew ground bidirectional
rlabel metal1 s -35 -3 -30 33 4 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 10 -3 15 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 28 -3 33 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 89 -3 94 25 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 145 -3 150 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 180 -3 185 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 225 -3 230 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s 260 -3 265 33 6 VSS
port 8 nsew ground bidirectional
rlabel metal1 s -81 -3 293 9 6 VSS
port 8 nsew ground bidirectional
<< properties >>
string FIXED_BBOX -81 -3 293 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
