magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 2248
<< mvpmos >>
rect 0 0 120 2128
rect 224 0 344 2128
<< mvpdiff >>
rect -88 2115 0 2128
rect -88 1661 -75 2115
rect -29 1661 0 2115
rect -88 1604 0 1661
rect -88 1558 -75 1604
rect -29 1558 0 1604
rect -88 1501 0 1558
rect -88 1455 -75 1501
rect -29 1455 0 1501
rect -88 1398 0 1455
rect -88 1352 -75 1398
rect -29 1352 0 1398
rect -88 1295 0 1352
rect -88 1249 -75 1295
rect -29 1249 0 1295
rect -88 1192 0 1249
rect -88 1146 -75 1192
rect -29 1146 0 1192
rect -88 1089 0 1146
rect -88 1043 -75 1089
rect -29 1043 0 1089
rect -88 986 0 1043
rect -88 940 -75 986
rect -29 940 0 986
rect -88 883 0 940
rect -88 837 -75 883
rect -29 837 0 883
rect -88 780 0 837
rect -88 734 -75 780
rect -29 734 0 780
rect -88 677 0 734
rect -88 631 -75 677
rect -29 631 0 677
rect -88 574 0 631
rect -88 528 -75 574
rect -29 528 0 574
rect -88 471 0 528
rect -88 425 -75 471
rect -29 425 0 471
rect -88 368 0 425
rect -88 322 -75 368
rect -29 322 0 368
rect -88 265 0 322
rect -88 219 -75 265
rect -29 219 0 265
rect -88 162 0 219
rect -88 116 -75 162
rect -29 116 0 162
rect -88 59 0 116
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 2115 224 2128
rect 120 1661 149 2115
rect 195 1661 224 2115
rect 120 1604 224 1661
rect 120 1558 149 1604
rect 195 1558 224 1604
rect 120 1501 224 1558
rect 120 1455 149 1501
rect 195 1455 224 1501
rect 120 1398 224 1455
rect 120 1352 149 1398
rect 195 1352 224 1398
rect 120 1295 224 1352
rect 120 1249 149 1295
rect 195 1249 224 1295
rect 120 1192 224 1249
rect 120 1146 149 1192
rect 195 1146 224 1192
rect 120 1089 224 1146
rect 120 1043 149 1089
rect 195 1043 224 1089
rect 120 986 224 1043
rect 120 940 149 986
rect 195 940 224 986
rect 120 883 224 940
rect 120 837 149 883
rect 195 837 224 883
rect 120 780 224 837
rect 120 734 149 780
rect 195 734 224 780
rect 120 677 224 734
rect 120 631 149 677
rect 195 631 224 677
rect 120 574 224 631
rect 120 528 149 574
rect 195 528 224 574
rect 120 471 224 528
rect 120 425 149 471
rect 195 425 224 471
rect 120 368 224 425
rect 120 322 149 368
rect 195 322 224 368
rect 120 265 224 322
rect 120 219 149 265
rect 195 219 224 265
rect 120 162 224 219
rect 120 116 149 162
rect 195 116 224 162
rect 120 59 224 116
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 2115 432 2128
rect 344 1661 373 2115
rect 419 1661 432 2115
rect 344 1604 432 1661
rect 344 1558 373 1604
rect 419 1558 432 1604
rect 344 1501 432 1558
rect 344 1455 373 1501
rect 419 1455 432 1501
rect 344 1398 432 1455
rect 344 1352 373 1398
rect 419 1352 432 1398
rect 344 1295 432 1352
rect 344 1249 373 1295
rect 419 1249 432 1295
rect 344 1192 432 1249
rect 344 1146 373 1192
rect 419 1146 432 1192
rect 344 1089 432 1146
rect 344 1043 373 1089
rect 419 1043 432 1089
rect 344 986 432 1043
rect 344 940 373 986
rect 419 940 432 986
rect 344 883 432 940
rect 344 837 373 883
rect 419 837 432 883
rect 344 780 432 837
rect 344 734 373 780
rect 419 734 432 780
rect 344 677 432 734
rect 344 631 373 677
rect 419 631 432 677
rect 344 574 432 631
rect 344 528 373 574
rect 419 528 432 574
rect 344 471 432 528
rect 344 425 373 471
rect 419 425 432 471
rect 344 368 432 425
rect 344 322 373 368
rect 419 322 432 368
rect 344 265 432 322
rect 344 219 373 265
rect 419 219 432 265
rect 344 162 432 219
rect 344 116 373 162
rect 419 116 432 162
rect 344 59 432 116
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 1661 -29 2115
rect -75 1558 -29 1604
rect -75 1455 -29 1501
rect -75 1352 -29 1398
rect -75 1249 -29 1295
rect -75 1146 -29 1192
rect -75 1043 -29 1089
rect -75 940 -29 986
rect -75 837 -29 883
rect -75 734 -29 780
rect -75 631 -29 677
rect -75 528 -29 574
rect -75 425 -29 471
rect -75 322 -29 368
rect -75 219 -29 265
rect -75 116 -29 162
rect -75 13 -29 59
rect 149 1661 195 2115
rect 149 1558 195 1604
rect 149 1455 195 1501
rect 149 1352 195 1398
rect 149 1249 195 1295
rect 149 1146 195 1192
rect 149 1043 195 1089
rect 149 940 195 986
rect 149 837 195 883
rect 149 734 195 780
rect 149 631 195 677
rect 149 528 195 574
rect 149 425 195 471
rect 149 322 195 368
rect 149 219 195 265
rect 149 116 195 162
rect 149 13 195 59
rect 373 1661 419 2115
rect 373 1558 419 1604
rect 373 1455 419 1501
rect 373 1352 419 1398
rect 373 1249 419 1295
rect 373 1146 419 1192
rect 373 1043 419 1089
rect 373 940 419 986
rect 373 837 419 883
rect 373 734 419 780
rect 373 631 419 677
rect 373 528 419 574
rect 373 425 419 471
rect 373 322 419 368
rect 373 219 419 265
rect 373 116 419 162
rect 373 13 419 59
<< polysilicon >>
rect 0 2128 120 2172
rect 224 2128 344 2172
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 2115 -29 2128
rect -75 1604 -29 1661
rect -75 1501 -29 1558
rect -75 1398 -29 1455
rect -75 1295 -29 1352
rect -75 1192 -29 1249
rect -75 1089 -29 1146
rect -75 986 -29 1043
rect -75 883 -29 940
rect -75 780 -29 837
rect -75 677 -29 734
rect -75 574 -29 631
rect -75 471 -29 528
rect -75 368 -29 425
rect -75 265 -29 322
rect -75 162 -29 219
rect -75 59 -29 116
rect -75 0 -29 13
rect 149 2115 195 2128
rect 149 1604 195 1661
rect 149 1501 195 1558
rect 149 1398 195 1455
rect 149 1295 195 1352
rect 149 1192 195 1249
rect 149 1089 195 1146
rect 149 986 195 1043
rect 149 883 195 940
rect 149 780 195 837
rect 149 677 195 734
rect 149 574 195 631
rect 149 471 195 528
rect 149 368 195 425
rect 149 265 195 322
rect 149 162 195 219
rect 149 59 195 116
rect 149 0 195 13
rect 373 2115 419 2128
rect 373 1604 419 1661
rect 373 1501 419 1558
rect 373 1398 419 1455
rect 373 1295 419 1352
rect 373 1192 419 1249
rect 373 1089 419 1146
rect 373 986 419 1043
rect 373 883 419 940
rect 373 780 419 837
rect 373 677 419 734
rect 373 574 419 631
rect 373 471 419 528
rect 373 368 419 425
rect 373 265 419 322
rect 373 162 419 219
rect 373 59 419 116
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 1064 -52 1064 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 1064 396 1064 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 1064 172 1064 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 707044
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 701670
<< end >>
