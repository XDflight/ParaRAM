magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 1342 23867 22665 29129
rect 1216 17407 22310 19961
rect 22338 17406 22926 19961
rect 22827 14326 23842 15917
rect 22880 8391 23005 9181
<< mvpmos >>
rect 6089 27950 6209 28632
rect 6314 27950 6434 28632
rect 6780 27950 6900 28632
rect 7005 27950 7125 28632
rect 16889 27950 17009 28632
rect 17114 27950 17234 28632
rect 17580 27950 17700 28632
rect 17805 27950 17925 28632
rect 6089 27175 6209 27857
rect 6314 27175 6434 27857
rect 6780 27175 6900 27857
rect 7005 27175 7125 27857
rect 16889 27175 17009 27857
rect 17114 27175 17234 27857
rect 17580 27175 17700 27857
rect 17805 27175 17925 27857
<< mvpdiff >>
rect 5983 27950 6089 28632
rect 6209 27950 6314 28632
rect 6434 27950 6540 28632
rect 6674 27950 6780 28632
rect 6900 27950 7005 28632
rect 7125 27950 7231 28632
rect 16783 27950 16889 28632
rect 17009 27950 17114 28632
rect 17234 27950 17340 28632
rect 17474 27950 17580 28632
rect 17700 27950 17805 28632
rect 17925 27950 18031 28632
rect 5983 27175 6089 27857
rect 6209 27175 6314 27857
rect 6434 27175 6540 27857
rect 6674 27175 6780 27857
rect 6900 27175 7005 27857
rect 7125 27175 7231 27857
rect 16783 27175 16889 27857
rect 17009 27175 17114 27857
rect 17234 27175 17340 27857
rect 17474 27175 17580 27857
rect 17700 27175 17805 27857
rect 17925 27175 18031 27857
<< metal1 >>
rect 936 29878 1116 29890
rect 936 29826 948 29878
rect 1104 29826 1116 29878
rect 936 29814 1116 29826
rect 1125 29774 1289 30213
rect 6525 29774 6689 30213
rect 11925 29890 12089 30213
rect 11777 29878 12089 29890
rect 11777 29826 11789 29878
rect 11945 29826 12089 29878
rect 11777 29814 12089 29826
rect 11925 29774 12089 29814
rect 17325 29774 17489 30213
rect 22725 29997 22889 30213
rect 22725 29985 22988 29997
rect 22725 29933 22800 29985
rect 22852 29933 22924 29985
rect 22976 29933 22988 29985
rect 22725 29890 22988 29933
rect 22559 29861 25315 29890
rect 22559 29809 22800 29861
rect 22852 29809 22924 29861
rect 22976 29809 25315 29861
rect 22559 29720 25315 29809
rect 22263 27031 22913 27105
rect 23206 18457 23552 19818
rect 23259 4973 23599 5013
rect 23259 4921 23297 4973
rect 23349 4921 23509 4973
rect 23561 4921 23599 4973
rect 23259 4755 23599 4921
rect 23259 4703 23297 4755
rect 23349 4703 23509 4755
rect 23561 4703 23599 4755
rect 23259 4662 23599 4703
<< via1 >>
rect 948 29826 1104 29878
rect 11789 29826 11945 29878
rect 22800 29933 22852 29985
rect 22924 29933 22976 29985
rect 22800 29809 22852 29861
rect 22924 29809 22976 29861
rect 23297 4921 23349 4973
rect 23509 4921 23561 4973
rect 23297 4703 23349 4755
rect 23509 4703 23561 4755
<< metal2 >>
rect 976 29987 1077 31182
rect 976 29931 996 29987
rect 1052 29931 1077 29987
rect 976 29890 1077 29931
rect 936 29878 1116 29890
rect 936 29826 948 29878
rect 1104 29826 1116 29878
rect 936 29814 996 29826
rect 976 29799 996 29814
rect 1052 29814 1116 29826
rect 1052 29799 1077 29814
rect 976 29723 1077 29799
rect 976 29667 996 29723
rect 1052 29667 1077 29723
rect 976 29591 1077 29667
rect 976 29535 996 29591
rect 1052 29535 1077 29591
rect 976 29471 1077 29535
rect 1337 27527 1437 31182
rect 11777 29987 11877 31182
rect 11777 29931 11798 29987
rect 11854 29931 11877 29987
rect 11777 29890 11877 29931
rect 11777 29878 11957 29890
rect 11777 29826 11789 29878
rect 11945 29826 11957 29878
rect 11777 29799 11798 29826
rect 11854 29814 11957 29826
rect 11854 29799 11877 29814
rect 11777 29723 11877 29799
rect 11777 29667 11798 29723
rect 11854 29667 11877 29723
rect 11777 29591 11877 29667
rect 11777 29535 11798 29591
rect 11854 29535 11877 29591
rect 11777 29471 11877 29535
rect 12137 27527 12237 31182
rect 22577 27527 22677 31182
rect 22937 29997 23037 31182
rect 22788 29987 23037 29997
rect 22788 29985 22958 29987
rect 22788 29933 22800 29985
rect 22852 29933 22924 29985
rect 22788 29931 22958 29933
rect 23014 29931 23037 29987
rect 22788 29861 23037 29931
rect 22788 29809 22800 29861
rect 22852 29809 22924 29861
rect 22976 29855 23037 29861
rect 22788 29799 22958 29809
rect 23014 29799 23037 29855
rect 22788 29797 23037 29799
rect 22937 29723 23037 29797
rect 22937 29667 22958 29723
rect 23014 29667 23037 29723
rect 22937 29591 23037 29667
rect 22937 29535 22958 29591
rect 23014 29535 23037 29591
rect 22937 27527 23037 29535
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4757 23599 4919
rect 23259 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 23259 4662 23599 4701
<< via2 >>
rect 996 29931 1052 29987
rect 996 29826 1052 29855
rect 996 29799 1052 29826
rect 996 29667 1052 29723
rect 996 29535 1052 29591
rect 11798 29931 11854 29987
rect 11798 29826 11854 29855
rect 11798 29799 11854 29826
rect 11798 29667 11854 29723
rect 11798 29535 11854 29591
rect 22958 29985 23014 29987
rect 22958 29933 22976 29985
rect 22976 29933 23014 29985
rect 22958 29931 23014 29933
rect 22958 29809 22976 29855
rect 22976 29809 23014 29855
rect 22958 29799 23014 29809
rect 22958 29667 23014 29723
rect 22958 29535 23014 29591
rect 23295 4973 23351 4975
rect 23295 4921 23297 4973
rect 23297 4921 23349 4973
rect 23349 4921 23351 4973
rect 23295 4919 23351 4921
rect 23507 4973 23563 4975
rect 23507 4921 23509 4973
rect 23509 4921 23561 4973
rect 23561 4921 23563 4973
rect 23507 4919 23563 4921
rect 23295 4755 23351 4757
rect 23295 4703 23297 4755
rect 23297 4703 23349 4755
rect 23349 4703 23351 4755
rect 23295 4701 23351 4703
rect 23507 4755 23563 4757
rect 23507 4703 23509 4755
rect 23509 4703 23561 4755
rect 23561 4703 23563 4755
rect 23507 4701 23563 4703
<< metal3 >>
rect -1 39107 23681 39307
rect -1 30537 23681 30897
rect 52 30139 23681 30279
rect 800 29987 24087 29997
rect 800 29943 996 29987
rect -1 29931 996 29943
rect 1052 29931 11798 29987
rect 11854 29931 22958 29987
rect 23014 29931 24087 29987
rect -1 29855 24087 29931
rect -1 29799 996 29855
rect 1052 29799 11798 29855
rect 11854 29799 22958 29855
rect 23014 29799 24087 29855
rect -1 29723 24087 29799
rect -1 29667 996 29723
rect 1052 29667 11798 29723
rect 11854 29667 22958 29723
rect 23014 29667 24087 29723
rect -1 29591 24087 29667
rect -1 29535 996 29591
rect 1052 29535 11798 29591
rect 11854 29535 22958 29591
rect 23014 29535 24087 29591
rect -1 29517 24087 29535
rect -1 29471 1243 29517
rect 800 27296 24087 29105
rect 1314 21089 23252 21304
rect 1314 20767 23252 20983
rect 1314 20446 23252 20661
rect 1314 20124 23252 20339
rect 1314 19432 23252 19648
rect 1314 19110 23252 19326
rect 1314 18789 23252 19004
rect 1314 18467 23252 18682
rect 1314 17918 23252 18361
rect 1314 16807 23252 17263
rect 1314 12996 23252 15720
rect 1314 9308 23252 12711
rect 1262 8442 23710 9158
rect 1262 7016 24488 7827
rect 1314 5154 23971 6474
rect 1165 4929 22567 5005
rect 23259 4975 23599 5014
rect 23259 4919 23295 4975
rect 23351 4919 23507 4975
rect 23563 4919 23599 4975
rect 23259 4758 23599 4919
rect 1165 4757 23599 4758
rect 1165 4701 23295 4757
rect 23351 4701 23507 4757
rect 23563 4701 23599 4757
rect 1165 4662 23599 4701
rect 1314 3133 24166 4495
rect 1314 1961 24276 2576
rect 1314 1286 23252 1855
rect 1314 747 24089 1179
rect 1314 155 24508 610
rect 1277 -959 24602 -504
rect 1277 -1599 23252 -1247
rect 1277 -2041 23252 -1953
rect 1277 -2517 23252 -2165
rect 1277 -3242 23252 -2787
use M2_M1$$43374636_64x8m81  M2_M1$$43374636_64x8m81_0
timestamp 1666464484
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_0
timestamp 1666464484
transform -1 0 11867 0 -1 29852
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_1
timestamp 1666464484
transform -1 0 1026 0 -1 29852
box 0 0 1 1
use M2_M14310589983225_64x8m81  M2_M14310589983225_64x8m81_0
timestamp 1666464484
transform -1 0 22888 0 -1 29897
box 0 0 1 1
use M3_M2$$201416748_64x8m81  M3_M2$$201416748_64x8m81_0
timestamp 1666464484
transform 1 0 23429 0 1 4838
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_0
timestamp 1666464484
transform 1 0 1024 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_1
timestamp 1666464484
transform 1 0 11826 0 1 29761
box 0 0 1 1
use M3_M24310589983226_64x8m81  M3_M24310589983226_64x8m81_2
timestamp 1666464484
transform 1 0 22986 0 1 29761
box 0 0 1 1
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_0
timestamp 1666464484
transform 1 0 12186 0 1 28317
box -38 -764 38 764
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_1
timestamp 1666464484
transform 1 0 22626 0 1 28317
box -38 -764 38 764
use M3_M24310589983227_64x8m81  M3_M24310589983227_64x8m81_2
timestamp 1666464484
transform 1 0 1386 0 1 28317
box -38 -764 38 764
use col_64a_64x8m81  col_64a_64x8m81_0
timestamp 1666464484
transform 1 0 907 0 1 31107
box -1997 -68 23144 7268
use dcap_103_novia_64x8m81  dcap_103_novia_64x8m81_0
array 0 35 619 0 0 0
timestamp 1666464484
transform 1 0 288 0 1 29009
box -203 -284 822 881
use rdummy_64x4_64x8m81  rdummy_64x4_64x8m81_0
timestamp 1666464484
transform 1 0 307 0 1 30207
box -269 -25410 24098 9088
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_0
timestamp 1666464484
transform -1 0 12194 0 1 6
box -269 -3400 7633 31133
use saout_R_m2_64x8m81  saout_R_m2_64x8m81_1
timestamp 1666464484
transform -1 0 22994 0 1 6
box -269 -3400 7633 31133
use saout_m2_64x8m81  saout_m2_64x8m81_0
timestamp 1666464484
transform 1 0 11820 0 1 -1
box -269 -3393 7633 31140
use saout_m2_64x8m81  saout_m2_64x8m81_1
timestamp 1666464484
transform 1 0 1020 0 1 -1
box -269 -3393 7633 31140
<< labels >>
rlabel metal1 s 7342 15928 7342 15928 4 pcb[6]
port 1 nsew
rlabel metal1 s 5921 15928 5921 15928 4 pcb[7]
port 2 nsew
rlabel metal1 s 18209 15928 18209 15928 4 pcb[4]
port 3 nsew
rlabel metal1 s 1827 18163 1827 18163 4 vdd
port 4 nsew
flabel metal1 s 22465 -3332 22465 -3332 0 FreeSans 600 0 0 0 WEN[4]
port 5 nsew
flabel metal1 s 1584 -3332 1584 -3332 0 FreeSans 600 0 0 0 WEN[7]
port 6 nsew
rlabel metal1 s 16588 15928 16588 15928 4 pcb[5]
port 7 nsew
flabel metal1 s 12358 -3332 12358 -3332 0 FreeSans 600 0 0 0 WEN[5]
port 8 nsew
flabel metal1 s 11643 -3332 11643 -3332 0 FreeSans 600 0 0 0 WEN[6]
port 9 nsew
rlabel metal3 s 1607 36968 1607 36968 4 WL[6]
port 10 nsew
rlabel metal3 s 1607 36068 1607 36068 4 WL[5]
port 11 nsew
rlabel metal3 s 1777 1467 1777 1467 4 men
port 12 nsew
rlabel metal3 s 1704 18914 1704 18914 4 ypass[1]
port 13 nsew
rlabel metal3 s 1704 19231 1704 19231 4 ypass[2]
port 14 nsew
rlabel metal3 s 1704 19548 1704 19548 4 ypass[3]
port 15 nsew
rlabel metal3 s 1704 20204 1704 20204 4 ypass[4]
port 16 nsew
rlabel metal3 s 1704 20528 1704 20528 4 ypass[5]
port 17 nsew
rlabel metal3 s 1704 20845 1704 20845 4 ypass[6]
port 18 nsew
rlabel metal3 s 1774 1467 1774 1467 4 men
port 12 nsew
rlabel metal3 s 1592 38757 1592 38757 4 DWL
port 19 nsew
rlabel metal3 s 1346 4726 1346 4726 4 tblhl
port 20 nsew
flabel metal3 s 1659 -2004 1659 -2004 0 FreeSans 1000 0 0 0 GWEN
port 21 nsew
flabel metal3 s 1659 -3019 1659 -3019 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
rlabel metal3 s 1777 8832 1777 8832 4 VDD
port 22 nsew
rlabel metal3 s 1777 5806 1777 5806 4 VSS
port 23 nsew
flabel metal3 s 1659 -781 1659 -781 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 -2347 1659 -2347 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
rlabel metal3 s 240 30277 240 30277 4 VSS
port 23 nsew
rlabel metal3 s 1777 39217 1777 39217 4 VSS
port 23 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 12 nsew
rlabel metal3 s 1704 18591 1704 18591 4 ypass[0]
port 24 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 12 nsew
rlabel metal3 s 1346 4983 1346 4983 4 GWE
port 25 nsew
rlabel metal3 s 1608 31568 1608 31568 4 WL[0]
port 26 nsew
rlabel metal3 s 1608 33368 1608 33368 4 WL[2]
port 27 nsew
rlabel metal3 s 1608 34268 1608 34268 4 WL[3]
port 28 nsew
rlabel metal3 s 1608 35168 1608 35168 4 WL[4]
port 29 nsew
rlabel metal3 s 1608 37868 1608 37868 4 WL[7]
port 30 nsew
rlabel metal3 s 1608 32468 1608 32468 4 WL[1]
port 31 nsew
rlabel metal3 s 1705 21162 1705 21162 4 ypass[7]
port 32 nsew
rlabel metal3 s 1777 1466 1777 1466 4 men
port 12 nsew
rlabel metal3 s 1775 1466 1775 1466 4 men
port 12 nsew
flabel metal3 s 1659 -1446 1659 -1446 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 390 1659 390 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 3623 1659 3623 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 7598 1659 7598 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 14001 1659 14001 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 18106 1659 18106 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 1659 28191 1659 28191 0 FreeSans 2000 0 0 0 VDD
port 22 nsew
flabel metal3 s 315 29699 315 29699 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 23123 1659 23123 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 16976 1659 16976 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 12236 1659 12236 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 6155 1659 6155 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 2247 1659 2247 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
flabel metal3 s 1659 949 1659 949 0 FreeSans 2000 0 0 0 VSS
port 23 nsew
rlabel metal2 s 1523 104 1523 104 4 din[4]
port 33 nsew
rlabel metal2 s 22489 104 22489 104 4 din[7]
port 34 nsew
rlabel metal2 s 10837 138 10837 138 4 q[5]
port 35 nsew
rlabel metal2 s 13166 104 13166 104 4 q[6]
port 36 nsew
rlabel metal2 s 21642 104 21642 104 4 q[7]
port 37 nsew
rlabel metal2 s 11684 104 11684 104 4 din[5]
port 38 nsew
rlabel metal2 s 12319 104 12319 104 4 din[6]
port 39 nsew
rlabel metal2 s 2377 104 2377 104 4 q[4]
port 40 nsew
<< properties >>
string GDS_END 2231038
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2220918
<< end >>
