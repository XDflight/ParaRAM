magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 424
rect 224 0 344 424
rect 448 0 568 424
rect 672 0 792 424
rect 896 0 1016 424
rect 1120 0 1240 424
<< mvndiff >>
rect -88 411 0 424
rect -88 365 -75 411
rect -29 365 0 411
rect -88 294 0 365
rect -88 248 -75 294
rect -29 248 0 294
rect -88 177 0 248
rect -88 131 -75 177
rect -29 131 0 177
rect -88 59 0 131
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 411 224 424
rect 120 365 149 411
rect 195 365 224 411
rect 120 294 224 365
rect 120 248 149 294
rect 195 248 224 294
rect 120 177 224 248
rect 120 131 149 177
rect 195 131 224 177
rect 120 59 224 131
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 411 448 424
rect 344 365 373 411
rect 419 365 448 411
rect 344 294 448 365
rect 344 248 373 294
rect 419 248 448 294
rect 344 177 448 248
rect 344 131 373 177
rect 419 131 448 177
rect 344 59 448 131
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 411 672 424
rect 568 365 597 411
rect 643 365 672 411
rect 568 294 672 365
rect 568 248 597 294
rect 643 248 672 294
rect 568 177 672 248
rect 568 131 597 177
rect 643 131 672 177
rect 568 59 672 131
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 411 896 424
rect 792 365 821 411
rect 867 365 896 411
rect 792 294 896 365
rect 792 248 821 294
rect 867 248 896 294
rect 792 177 896 248
rect 792 131 821 177
rect 867 131 896 177
rect 792 59 896 131
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 411 1120 424
rect 1016 365 1045 411
rect 1091 365 1120 411
rect 1016 294 1120 365
rect 1016 248 1045 294
rect 1091 248 1120 294
rect 1016 177 1120 248
rect 1016 131 1045 177
rect 1091 131 1120 177
rect 1016 59 1120 131
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 411 1328 424
rect 1240 365 1269 411
rect 1315 365 1328 411
rect 1240 294 1328 365
rect 1240 248 1269 294
rect 1315 248 1328 294
rect 1240 177 1328 248
rect 1240 131 1269 177
rect 1315 131 1328 177
rect 1240 59 1328 131
rect 1240 13 1269 59
rect 1315 13 1328 59
rect 1240 0 1328 13
<< mvndiffc >>
rect -75 365 -29 411
rect -75 248 -29 294
rect -75 131 -29 177
rect -75 13 -29 59
rect 149 365 195 411
rect 149 248 195 294
rect 149 131 195 177
rect 149 13 195 59
rect 373 365 419 411
rect 373 248 419 294
rect 373 131 419 177
rect 373 13 419 59
rect 597 365 643 411
rect 597 248 643 294
rect 597 131 643 177
rect 597 13 643 59
rect 821 365 867 411
rect 821 248 867 294
rect 821 131 867 177
rect 821 13 867 59
rect 1045 365 1091 411
rect 1045 248 1091 294
rect 1045 131 1091 177
rect 1045 13 1091 59
rect 1269 365 1315 411
rect 1269 248 1315 294
rect 1269 131 1315 177
rect 1269 13 1315 59
<< polysilicon >>
rect 0 424 120 468
rect 224 424 344 468
rect 448 424 568 468
rect 672 424 792 468
rect 896 424 1016 468
rect 1120 424 1240 468
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
<< metal1 >>
rect -75 411 -29 424
rect -75 294 -29 365
rect -75 177 -29 248
rect -75 59 -29 131
rect -75 0 -29 13
rect 149 411 195 424
rect 149 294 195 365
rect 149 177 195 248
rect 149 59 195 131
rect 149 0 195 13
rect 373 411 419 424
rect 373 294 419 365
rect 373 177 419 248
rect 373 59 419 131
rect 373 0 419 13
rect 597 411 643 424
rect 597 294 643 365
rect 597 177 643 248
rect 597 59 643 131
rect 597 0 643 13
rect 821 411 867 424
rect 821 294 867 365
rect 821 177 867 248
rect 821 59 867 131
rect 821 0 867 13
rect 1045 411 1091 424
rect 1045 294 1091 365
rect 1045 177 1091 248
rect 1045 59 1091 131
rect 1045 0 1091 13
rect 1269 411 1315 424
rect 1269 294 1315 365
rect 1269 177 1315 248
rect 1269 59 1315 131
rect 1269 0 1315 13
<< labels >>
flabel metal1 s -52 212 -52 212 0 FreeSans 200 0 0 0 S
flabel metal1 s 1292 212 1292 212 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 212 172 212 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 212 396 212 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 212 620 212 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 212 844 212 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 212 1068 212 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 365464
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 360866
<< end >>
