magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 272
<< mvndiff >>
rect -88 259 0 272
rect -88 13 -75 259
rect -29 13 0 259
rect -88 0 0 13
rect 120 259 208 272
rect 120 13 149 259
rect 195 13 208 259
rect 120 0 208 13
<< mvndiffc >>
rect -75 13 -29 259
rect 149 13 195 259
<< polysilicon >>
rect 0 272 120 316
rect 0 -44 120 0
<< metal1 >>
rect -75 259 -29 272
rect -75 0 -29 13
rect 149 259 195 272
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 136 -52 136 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 136 172 136 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 216302
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 215022
<< end >>
