magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 896 844
rect 281 602 349 724
rect 535 540 581 678
rect 728 602 796 724
rect 141 325 330 430
rect 535 442 760 540
rect 141 122 203 325
rect 696 260 760 442
rect 535 213 760 260
rect 281 60 349 153
rect 535 114 581 213
rect 748 60 816 153
rect 0 -60 896 60
<< obsm1 >>
rect 49 525 95 678
rect 49 478 426 525
rect 49 114 95 478
rect 380 378 426 478
rect 380 310 648 378
<< labels >>
rlabel metal1 s 141 325 330 430 6 I
port 1 nsew default input
rlabel metal1 s 141 122 203 325 6 I
port 1 nsew default input
rlabel metal1 s 535 540 581 678 6 Z
port 2 nsew default output
rlabel metal1 s 535 442 760 540 6 Z
port 2 nsew default output
rlabel metal1 s 696 260 760 442 6 Z
port 2 nsew default output
rlabel metal1 s 535 213 760 260 6 Z
port 2 nsew default output
rlabel metal1 s 535 114 581 213 6 Z
port 2 nsew default output
rlabel metal1 s 0 724 896 844 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 728 602 796 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 281 602 349 724 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 748 60 816 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 281 60 349 153 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 896 60 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1309198
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1306330
<< end >>
