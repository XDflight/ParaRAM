magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 243 595
<< polysilicon >>
rect -31 454 88 527
rect -31 -74 88 0
use pmos_5p04310589983214_64x8m81  pmos_5p04310589983214_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 574
<< properties >>
string GDS_END 263262
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 262948
<< end >>
