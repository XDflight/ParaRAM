magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 918 4480 1098
rect 294 685 340 918
rect 642 719 688 918
rect 1538 896 1584 918
rect 2166 896 2212 918
rect 2955 792 3023 918
rect 3363 792 3431 918
rect 3782 781 3828 918
rect 3930 775 3976 918
rect 4338 775 4384 918
rect 142 354 316 430
rect 678 354 866 430
rect 283 90 351 209
rect 688 90 734 285
rect 798 242 866 354
rect 1775 90 1843 274
rect 3054 242 3122 412
rect 3351 464 3554 542
rect 3374 90 3420 245
rect 3910 90 3956 233
rect 4134 169 4226 766
rect 4358 90 4404 233
rect 0 -90 4480 90
<< obsm1 >>
rect 90 621 136 737
rect 734 850 1195 868
rect 2491 850 2559 870
rect 734 804 2559 850
rect 734 643 780 804
rect 90 575 428 621
rect 382 308 428 575
rect 70 262 428 308
rect 498 597 780 643
rect 846 637 892 753
rect 70 238 116 262
rect 498 238 564 597
rect 846 591 958 637
rect 912 263 958 591
rect 1050 550 1096 753
rect 1304 690 1832 758
rect 1304 596 1350 690
rect 1930 661 1976 758
rect 1930 615 2156 661
rect 1930 596 1976 615
rect 2018 550 2064 569
rect 1050 504 2064 550
rect 1136 263 1182 504
rect 2018 501 2064 504
rect 2110 491 2156 615
rect 2414 491 2460 755
rect 1420 455 2001 458
rect 2110 455 2460 491
rect 1420 445 2460 455
rect 2618 746 2927 755
rect 2618 709 3738 746
rect 1272 344 1318 423
rect 1420 412 2288 445
rect 1420 390 1466 412
rect 1984 409 2288 412
rect 1506 344 1967 366
rect 1272 320 1967 344
rect 1272 298 1546 320
rect 1921 182 1967 320
rect 2242 263 2288 409
rect 2618 380 2664 709
rect 2899 700 3738 709
rect 2466 334 2664 380
rect 2466 263 2512 334
rect 2822 296 2868 661
rect 2690 274 2868 296
rect 2690 228 3008 274
rect 2962 196 3008 228
rect 3170 196 3216 645
rect 3578 582 3646 650
rect 3600 423 3646 582
rect 3692 485 3738 700
rect 3600 418 4064 423
rect 3275 372 4064 418
rect 3766 355 4064 372
rect 3766 263 3812 355
rect 1921 136 2876 182
rect 2962 150 3216 196
<< labels >>
rlabel metal1 s 678 354 866 430 6 D
port 1 nsew default input
rlabel metal1 s 798 242 866 354 6 D
port 1 nsew default input
rlabel metal1 s 3351 464 3554 542 6 RN
port 2 nsew default input
rlabel metal1 s 3054 242 3122 412 6 SETN
port 3 nsew default input
rlabel metal1 s 142 354 316 430 6 CLKN
port 4 nsew clock input
rlabel metal1 s 4134 169 4226 766 6 Q
port 5 nsew default output
rlabel metal1 s 0 918 4480 1098 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 896 4384 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 896 3976 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 896 3828 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3363 896 3431 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2955 896 3023 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2166 896 2212 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1538 896 1584 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 896 688 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 896 340 918 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 792 4384 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 792 3976 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 792 3828 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3363 792 3431 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2955 792 3023 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 792 688 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 792 340 896 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 781 4384 792 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 781 3976 792 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3782 781 3828 792 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 781 688 792 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 781 340 792 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 4338 775 4384 781 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3930 775 3976 781 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 775 688 781 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 775 340 781 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 642 719 688 775 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 719 340 775 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 294 685 340 719 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 688 274 734 285 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1775 245 1843 274 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 688 245 734 274 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3374 233 3420 245 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1775 233 1843 245 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 688 233 734 245 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4358 209 4404 233 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3910 209 3956 233 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3374 209 3420 233 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1775 209 1843 233 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 688 209 734 233 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 4358 90 4404 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3910 90 3956 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3374 90 3420 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1775 90 1843 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 688 90 734 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 283 90 351 209 6 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4480 90 8 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4480 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 530788
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 520688
<< end >>
