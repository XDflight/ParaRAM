magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< ndiff >>
rect -700 23 700 42
rect -700 -23 -681 23
rect 681 -23 700 23
rect -700 -42 700 -23
<< ndiffc >>
rect -681 -23 681 23
<< metal1 >>
rect -692 23 692 34
rect -692 -23 -681 23
rect 681 -23 692 23
rect -692 -34 692 -23
<< properties >>
string GDS_END 281118
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 279962
<< end >>
