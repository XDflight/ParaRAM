magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 7178 9364 8480 10100
rect 6657 6921 12228 7706
rect 6734 4159 12228 6921
rect 7398 1986 8542 1987
rect 9089 1986 10232 1987
rect 10779 1986 11923 1987
rect 6914 797 11923 1986
<< pmos >>
rect 7433 9505 7553 9960
rect 7657 9505 7777 9960
rect 7881 9505 8001 9960
rect 8105 9505 8225 9960
<< pdiff >>
rect 7314 9801 7433 9960
rect 7314 9755 7358 9801
rect 7404 9755 7433 9801
rect 7314 9597 7433 9755
rect 7314 9551 7358 9597
rect 7404 9551 7433 9597
rect 7314 9505 7433 9551
rect 7553 9505 7657 9960
rect 7777 9801 7881 9960
rect 7777 9755 7806 9801
rect 7852 9755 7881 9801
rect 7777 9597 7881 9755
rect 7777 9551 7806 9597
rect 7852 9551 7881 9597
rect 7777 9505 7881 9551
rect 8001 9505 8105 9960
rect 8225 9801 8344 9960
rect 8225 9755 8254 9801
rect 8300 9755 8344 9801
rect 8225 9597 8344 9755
rect 8225 9551 8254 9597
rect 8300 9551 8344 9597
rect 8225 9505 8344 9551
<< pdiffc >>
rect 7358 9755 7404 9801
rect 7358 9551 7404 9597
rect 7806 9755 7852 9801
rect 7806 9551 7852 9597
rect 8254 9755 8300 9801
rect 8254 9551 8300 9597
<< psubdiff >>
rect 8157 10830 12086 10889
rect 8157 10784 8287 10830
rect 8333 10784 8445 10830
rect 8491 10784 8603 10830
rect 8649 10784 8761 10830
rect 8807 10784 8919 10830
rect 8965 10784 9077 10830
rect 9123 10784 9235 10830
rect 9281 10784 9394 10830
rect 9440 10784 9552 10830
rect 9598 10784 9710 10830
rect 9756 10784 9868 10830
rect 9914 10784 10026 10830
rect 10072 10784 10184 10830
rect 10230 10784 10342 10830
rect 10388 10784 10500 10830
rect 10546 10784 10658 10830
rect 10704 10784 10817 10830
rect 10863 10784 10975 10830
rect 11021 10784 11133 10830
rect 11179 10784 11291 10830
rect 11337 10784 11449 10830
rect 11495 10784 11607 10830
rect 11653 10784 11765 10830
rect 11811 10784 11923 10830
rect 11969 10784 12086 10830
rect 8157 10724 12086 10784
<< psubdiffcont >>
rect 8287 10784 8333 10830
rect 8445 10784 8491 10830
rect 8603 10784 8649 10830
rect 8761 10784 8807 10830
rect 8919 10784 8965 10830
rect 9077 10784 9123 10830
rect 9235 10784 9281 10830
rect 9394 10784 9440 10830
rect 9552 10784 9598 10830
rect 9710 10784 9756 10830
rect 9868 10784 9914 10830
rect 10026 10784 10072 10830
rect 10184 10784 10230 10830
rect 10342 10784 10388 10830
rect 10500 10784 10546 10830
rect 10658 10784 10704 10830
rect 10817 10784 10863 10830
rect 10975 10784 11021 10830
rect 11133 10784 11179 10830
rect 11291 10784 11337 10830
rect 11449 10784 11495 10830
rect 11607 10784 11653 10830
rect 11765 10784 11811 10830
rect 11923 10784 11969 10830
<< polysilicon >>
rect 7965 10456 8049 10475
rect 7965 10316 7984 10456
rect 8030 10316 8049 10456
rect 7433 10159 7553 10209
rect 7148 10113 7553 10159
rect 7148 10067 7222 10113
rect 7268 10067 7380 10113
rect 7426 10067 7553 10113
rect 7148 10021 7553 10067
rect 7433 9960 7553 10021
rect 7657 10180 7777 10209
rect 7965 10180 8049 10316
rect 7657 10117 8049 10180
rect 7657 10095 8001 10117
rect 7657 9960 7777 10095
rect 7881 9960 8001 10095
rect 8105 10085 8309 10104
rect 8105 10039 8244 10085
rect 8290 10039 8309 10085
rect 8105 10020 8309 10039
rect 8105 9960 8225 10020
rect 9028 9996 9148 10205
rect 8909 9921 9253 9996
rect 7433 9432 7553 9505
rect 7657 9432 7777 9505
rect 7881 9432 8001 9505
rect 8105 9432 8225 9505
rect 8909 9459 9029 9921
rect 9133 9459 9253 9921
rect 8909 9440 9253 9459
rect 8909 9394 8953 9440
rect 9187 9394 9253 9440
rect 8909 9375 9253 9394
rect 303 4183 496 4228
rect 303 4137 377 4183
rect 423 4137 496 4183
rect 303 4091 496 4137
rect 1423 4183 1616 4228
rect 1423 4137 1497 4183
rect 1543 4137 1616 4183
rect 1423 4091 1616 4137
rect 1936 4183 2129 4228
rect 1936 4137 2010 4183
rect 2056 4137 2129 4183
rect 1936 4091 2129 4137
rect 3056 4183 3249 4228
rect 3056 4137 3130 4183
rect 3176 4137 3249 4183
rect 3056 4091 3249 4137
rect 527 3983 720 4028
rect 527 3937 601 3983
rect 647 3937 720 3983
rect 527 3891 720 3937
rect 1199 3983 1392 4028
rect 1199 3937 1273 3983
rect 1319 3937 1392 3983
rect 1199 3891 1392 3937
rect 3794 3983 3987 4028
rect 3794 3937 3868 3983
rect 3914 3937 3987 3983
rect 3794 3891 3987 3937
rect 4466 3983 4659 4028
rect 4466 3937 4540 3983
rect 4586 3937 4659 3983
rect 4466 3891 4659 3937
rect 751 3779 944 3824
rect 751 3733 825 3779
rect 871 3733 944 3779
rect 751 3687 944 3733
rect 2384 3779 2577 3824
rect 2384 3733 2458 3779
rect 2504 3733 2577 3779
rect 2384 3687 2577 3733
rect 4018 3779 4211 3824
rect 4018 3733 4092 3779
rect 4138 3733 4211 3779
rect 4018 3687 4211 3733
rect 5652 3779 5845 3824
rect 5652 3733 5726 3779
rect 5772 3733 5845 3779
rect 5652 3687 5845 3733
rect 3570 3578 3763 3623
rect 3570 3532 3644 3578
rect 3690 3532 3763 3578
rect 3570 3486 3763 3532
rect 4690 3578 4883 3623
rect 4690 3532 4764 3578
rect 4810 3532 4883 3578
rect 4690 3486 4883 3532
rect 5204 3578 5397 3623
rect 5204 3532 5278 3578
rect 5324 3532 5397 3578
rect 5204 3486 5397 3532
rect 6324 3578 6517 3623
rect 6324 3532 6398 3578
rect 6444 3532 6517 3578
rect 6324 3486 6517 3532
rect 2160 3376 2353 3421
rect 2160 3330 2234 3376
rect 2280 3330 2353 3376
rect 2160 3284 2353 3330
rect 2832 3376 3025 3421
rect 2832 3330 2906 3376
rect 2952 3330 3025 3376
rect 2832 3284 3025 3330
rect 5428 3376 5621 3421
rect 5428 3330 5502 3376
rect 5548 3330 5621 3376
rect 5428 3284 5621 3330
rect 6100 3376 6293 3421
rect 6100 3330 6174 3376
rect 6220 3330 6293 3376
rect 6100 3284 6293 3330
rect 975 3174 1168 3219
rect 975 3128 1049 3174
rect 1095 3128 1168 3174
rect 975 3082 1168 3128
rect 2608 3174 2801 3219
rect 2608 3128 2682 3174
rect 2728 3128 2801 3174
rect 2608 3082 2801 3128
rect 4242 3174 4435 3219
rect 4242 3128 4316 3174
rect 4362 3128 4435 3174
rect 4242 3082 4435 3128
rect 5876 3174 6069 3219
rect 5876 3128 5950 3174
rect 5996 3128 6069 3174
rect 5876 3082 6069 3128
<< polycontact >>
rect 7984 10316 8030 10456
rect 7222 10067 7268 10113
rect 7380 10067 7426 10113
rect 8244 10039 8290 10085
rect 8953 9394 9187 9440
rect 377 4137 423 4183
rect 1497 4137 1543 4183
rect 2010 4137 2056 4183
rect 3130 4137 3176 4183
rect 601 3937 647 3983
rect 1273 3937 1319 3983
rect 3868 3937 3914 3983
rect 4540 3937 4586 3983
rect 825 3733 871 3779
rect 2458 3733 2504 3779
rect 4092 3733 4138 3779
rect 5726 3733 5772 3779
rect 3644 3532 3690 3578
rect 4764 3532 4810 3578
rect 5278 3532 5324 3578
rect 6398 3532 6444 3578
rect 2234 3330 2280 3376
rect 2906 3330 2952 3376
rect 5502 3330 5548 3376
rect 6174 3330 6220 3376
rect 1049 3128 1095 3174
rect 2682 3128 2728 3174
rect 4316 3128 4362 3174
rect 5950 3128 5996 3174
<< metal1 >>
rect 6622 10830 12086 10880
rect 6622 10820 8287 10830
rect 6622 10768 7348 10820
rect 7400 10768 7787 10820
rect 7839 10784 8287 10820
rect 8333 10784 8445 10830
rect 8491 10784 8603 10830
rect 8649 10784 8761 10830
rect 8807 10784 8919 10830
rect 8965 10784 9077 10830
rect 9123 10784 9235 10830
rect 9281 10784 9394 10830
rect 9440 10784 9552 10830
rect 9598 10784 9710 10830
rect 9756 10784 9868 10830
rect 9914 10784 10026 10830
rect 10072 10784 10184 10830
rect 10230 10784 10342 10830
rect 10388 10784 10500 10830
rect 10546 10784 10658 10830
rect 10704 10784 10817 10830
rect 10863 10784 10975 10830
rect 11021 10784 11133 10830
rect 11179 10784 11291 10830
rect 11337 10784 11449 10830
rect 11495 10784 11607 10830
rect 11653 10784 11765 10830
rect 11811 10784 11923 10830
rect 11969 10784 12086 10830
rect 7839 10768 12086 10784
rect 6622 10763 12086 10768
rect 6622 10733 9171 10763
rect 7310 10602 7439 10733
rect 7310 10550 7348 10602
rect 7400 10550 7439 10602
rect 7749 10602 7887 10733
rect 9133 10711 9171 10733
rect 9223 10733 12086 10763
rect 9223 10711 9261 10733
rect 7310 10384 7439 10550
rect 7310 10332 7348 10384
rect 7400 10332 7439 10384
rect 7310 10292 7439 10332
rect 7323 10248 7439 10292
rect 7121 10114 7461 10155
rect 7121 10062 7159 10114
rect 7211 10113 7371 10114
rect 7423 10113 7461 10114
rect 7211 10067 7222 10113
rect 7268 10067 7371 10113
rect 7426 10067 7461 10113
rect 7211 10062 7371 10067
rect 7423 10062 7461 10067
rect 7121 10022 7461 10062
rect 7547 10152 7663 10554
rect 7749 10550 7787 10602
rect 7839 10550 7887 10602
rect 7749 10384 7887 10550
rect 7749 10332 7787 10384
rect 7839 10332 7887 10384
rect 7749 10292 7887 10332
rect 7971 10604 8095 10644
rect 7971 10552 8007 10604
rect 8059 10552 8095 10604
rect 7971 10456 8095 10552
rect 7971 10316 7984 10456
rect 8030 10386 8095 10456
rect 9133 10545 9261 10711
rect 9133 10493 9171 10545
rect 9223 10493 9261 10545
rect 8059 10334 8095 10386
rect 8030 10316 8095 10334
rect 7971 10294 8095 10316
rect 7771 10248 7887 10292
rect 7547 10033 7887 10152
rect 8917 10111 9033 10418
rect 9133 10327 9261 10493
rect 9133 10275 9171 10327
rect 9223 10275 9261 10327
rect 9133 10235 9261 10275
rect 10167 10112 10291 10145
rect 10165 10111 10294 10112
rect 8917 10105 10294 10111
rect 7323 9837 7439 9919
rect 7312 9801 7439 9837
rect 7312 9797 7358 9801
rect 7312 9745 7348 9797
rect 7404 9755 7439 9801
rect 7400 9745 7439 9755
rect 7312 9597 7439 9745
rect 7312 9579 7358 9597
rect 7312 9527 7348 9579
rect 7404 9551 7439 9597
rect 7400 9527 7439 9551
rect 7312 9514 7439 9527
rect 7771 9801 7887 10033
rect 8121 10092 8301 10104
rect 8121 10040 8133 10092
rect 8289 10085 8301 10092
rect 8121 10039 8244 10040
rect 8290 10039 8301 10085
rect 8121 10028 8301 10039
rect 8917 10053 10203 10105
rect 10255 10053 10294 10105
rect 8917 9978 10294 10053
rect 7771 9755 7806 9801
rect 7852 9755 7887 9801
rect 7771 9597 7887 9755
rect 7771 9551 7806 9597
rect 7852 9551 7887 9597
rect 7312 9487 7436 9514
rect 7771 9434 7887 9551
rect 8219 9851 8335 9919
rect 8498 9856 8622 9896
rect 8498 9851 8534 9856
rect 8219 9804 8534 9851
rect 8586 9851 8622 9856
rect 8586 9804 8915 9851
rect 8219 9801 8915 9804
rect 8219 9755 8254 9801
rect 8300 9755 8915 9801
rect 8219 9638 8915 9755
rect 8219 9597 8534 9638
rect 8219 9551 8254 9597
rect 8300 9586 8534 9597
rect 8586 9586 8915 9638
rect 9023 9616 9139 9978
rect 10167 9887 10291 9978
rect 9247 9811 9652 9851
rect 9247 9759 9562 9811
rect 9614 9759 9652 9811
rect 10167 9835 10203 9887
rect 10255 9835 10291 9887
rect 10167 9795 10291 9835
rect 8300 9551 8915 9586
rect 8219 9527 8915 9551
rect 9247 9593 9652 9759
rect 9247 9541 9562 9593
rect 9614 9541 9652 9593
rect 9247 9527 9652 9541
rect 8219 9514 8335 9527
rect 9526 9501 9650 9527
rect 8942 9440 9198 9451
rect 8942 9434 8953 9440
rect 7771 9394 8953 9434
rect 9187 9394 9198 9440
rect 7771 9393 9198 9394
rect 7771 9341 8430 9393
rect 8482 9341 8642 9393
rect 8694 9341 9198 9393
rect 7771 9314 9198 9341
rect 8392 9301 8732 9314
rect 7705 4659 7821 4660
rect 342 4183 457 4219
rect 342 4137 377 4183
rect 423 4137 457 4183
rect 342 4100 457 4137
rect 1462 4183 1577 4219
rect 1462 4137 1497 4183
rect 1543 4137 1577 4183
rect 1462 4100 1577 4137
rect 1975 4183 2090 4219
rect 1975 4137 2010 4183
rect 2056 4137 2090 4183
rect 1975 4100 2090 4137
rect 3095 4183 3210 4219
rect 3095 4137 3130 4183
rect 3176 4137 3210 4183
rect 3095 4100 3210 4137
rect 7698 4114 7828 4659
rect 566 3983 681 4019
rect 566 3937 601 3983
rect 647 3937 681 3983
rect 566 3900 681 3937
rect 1238 3983 1353 4019
rect 1238 3937 1273 3983
rect 1319 3937 1353 3983
rect 1238 3900 1353 3937
rect 3833 3983 3948 4019
rect 3833 3937 3868 3983
rect 3914 3937 3948 3983
rect 3833 3900 3948 3937
rect 4505 3983 4620 4019
rect 4505 3937 4540 3983
rect 4586 3937 4620 3983
rect 4505 3900 4620 3937
rect 9389 3984 9518 4025
rect 9389 3932 9428 3984
rect 9480 3932 9518 3984
rect 9389 3891 9518 3932
rect 790 3779 905 3815
rect 790 3733 825 3779
rect 871 3733 905 3779
rect 790 3696 905 3733
rect 2423 3779 2538 3815
rect 2423 3733 2458 3779
rect 2504 3733 2538 3779
rect 2423 3696 2538 3733
rect 4057 3779 4172 3815
rect 4057 3733 4092 3779
rect 4138 3733 4172 3779
rect 4057 3696 4172 3733
rect 5691 3779 5806 3815
rect 5691 3733 5726 3779
rect 5772 3733 5806 3779
rect 5691 3696 5806 3733
rect 11080 3782 11209 3823
rect 11080 3730 11119 3782
rect 11171 3730 11209 3782
rect 11080 3689 11209 3730
rect 3609 3578 3724 3614
rect 3609 3532 3644 3578
rect 3690 3532 3724 3578
rect 3609 3495 3724 3532
rect 4729 3578 4844 3614
rect 4729 3532 4764 3578
rect 4810 3532 4844 3578
rect 4729 3495 4844 3532
rect 5243 3578 5358 3614
rect 5243 3532 5278 3578
rect 5324 3532 5358 3578
rect 5243 3495 5358 3532
rect 6363 3578 6478 3614
rect 6363 3532 6398 3578
rect 6444 3532 6478 3578
rect 6363 3495 6478 3532
rect 8212 3581 8341 3622
rect 8212 3529 8251 3581
rect 8303 3529 8341 3581
rect 8212 3488 8341 3529
rect 2199 3376 2314 3412
rect 2199 3330 2234 3376
rect 2280 3330 2314 3376
rect 2199 3293 2314 3330
rect 2871 3376 2986 3412
rect 2871 3330 2906 3376
rect 2952 3330 2986 3376
rect 2871 3293 2986 3330
rect 5467 3376 5582 3412
rect 5467 3330 5502 3376
rect 5548 3330 5582 3376
rect 5467 3293 5582 3330
rect 6139 3376 6254 3412
rect 6139 3330 6174 3376
rect 6220 3330 6254 3376
rect 6139 3293 6254 3330
rect 9903 3379 10032 3420
rect 9903 3327 9942 3379
rect 9994 3327 10032 3379
rect 9903 3286 10032 3327
rect 1014 3174 1129 3210
rect 1014 3128 1049 3174
rect 1095 3128 1129 3174
rect 1014 3091 1129 3128
rect 2647 3174 2762 3210
rect 2647 3128 2682 3174
rect 2728 3128 2762 3174
rect 2647 3091 2762 3128
rect 4281 3174 4396 3210
rect 4281 3128 4316 3174
rect 4362 3128 4396 3174
rect 4281 3091 4396 3128
rect 5915 3174 6030 3210
rect 5915 3128 5950 3174
rect 5996 3128 6030 3174
rect 5915 3091 6030 3128
rect 11594 3177 11723 3218
rect 11594 3125 11633 3177
rect 11685 3125 11723 3177
rect 11594 3084 11723 3125
<< via1 >>
rect 7348 10768 7400 10820
rect 7787 10768 7839 10820
rect 7348 10550 7400 10602
rect 9171 10711 9223 10763
rect 7348 10332 7400 10384
rect 7159 10062 7211 10114
rect 7371 10113 7423 10114
rect 7371 10067 7380 10113
rect 7380 10067 7423 10113
rect 7371 10062 7423 10067
rect 7787 10550 7839 10602
rect 7787 10332 7839 10384
rect 8007 10552 8059 10604
rect 9171 10493 9223 10545
rect 8007 10334 8030 10386
rect 8030 10334 8059 10386
rect 9171 10275 9223 10327
rect 7348 9755 7358 9797
rect 7358 9755 7400 9797
rect 7348 9745 7400 9755
rect 7348 9551 7358 9579
rect 7358 9551 7400 9579
rect 7348 9527 7400 9551
rect 8133 10085 8289 10092
rect 8133 10040 8244 10085
rect 8244 10040 8289 10085
rect 10203 10053 10255 10105
rect 8534 9804 8586 9856
rect 8534 9586 8586 9638
rect 9562 9759 9614 9811
rect 10203 9835 10255 9887
rect 9562 9541 9614 9593
rect 8430 9341 8482 9393
rect 8642 9341 8694 9393
rect 9428 3932 9480 3984
rect 11119 3730 11171 3782
rect 8251 3529 8303 3581
rect 9942 3327 9994 3379
rect 11633 3125 11685 3177
<< metal2 >>
rect 719 10838 849 10971
rect 1073 10838 1202 10971
rect 2353 10838 2482 10971
rect 2715 10838 2845 10971
rect 3985 10838 4114 10971
rect 4338 10838 4468 10971
rect 5645 10838 5774 10971
rect 5968 10838 6097 10971
rect 7310 10822 7438 10859
rect 7310 10766 7346 10822
rect 7402 10766 7438 10822
rect 7310 10604 7438 10766
rect 7310 10548 7346 10604
rect 7402 10548 7438 10604
rect 7310 10386 7438 10548
rect 7310 10330 7346 10386
rect 7402 10330 7438 10386
rect 7310 10292 7438 10330
rect 7749 10822 7877 10859
rect 7749 10766 7785 10822
rect 7841 10766 7877 10822
rect 7749 10604 7877 10766
rect 9133 10765 9261 10802
rect 9133 10709 9169 10765
rect 9225 10709 9261 10765
rect 7749 10548 7785 10604
rect 7841 10548 7877 10604
rect 7749 10386 7877 10548
rect 7969 10604 8098 10645
rect 7969 10552 8007 10604
rect 8059 10552 8098 10604
rect 7969 10511 8098 10552
rect 9133 10547 9261 10709
rect 7749 10330 7785 10386
rect 7841 10330 7877 10386
rect 7749 10292 7877 10330
rect 7971 10386 8095 10511
rect 7971 10334 8007 10386
rect 8059 10334 8095 10386
rect 7971 10294 8095 10334
rect 9133 10491 9169 10547
rect 9225 10491 9261 10547
rect 9133 10329 9261 10491
rect 9133 10273 9169 10329
rect 9225 10273 9261 10329
rect 9133 10235 9261 10273
rect 7121 10114 8352 10155
rect 7121 10062 7159 10114
rect 7211 10062 7371 10114
rect 7423 10092 8352 10114
rect 7423 10062 8133 10092
rect 7121 10040 8133 10062
rect 8289 10040 8352 10092
rect 7121 10021 8352 10040
rect 10167 10105 10291 10145
rect 10167 10053 10203 10105
rect 10255 10053 10291 10105
rect 10167 9964 10291 10053
rect 8497 9858 8622 9897
rect 7311 9799 7436 9838
rect 7311 9743 7346 9799
rect 7402 9743 7436 9799
rect 7311 9581 7436 9743
rect 7311 9525 7346 9581
rect 7402 9525 7436 9581
rect 8497 9802 8532 9858
rect 8588 9802 8622 9858
rect 10165 9887 10294 9964
rect 8497 9640 8622 9802
rect 8497 9584 8532 9640
rect 8588 9584 8622 9640
rect 8497 9546 8622 9584
rect 9525 9813 9650 9852
rect 9525 9757 9560 9813
rect 9616 9757 9650 9813
rect 9525 9595 9650 9757
rect 7311 9487 7436 9525
rect 9525 9539 9560 9595
rect 9616 9539 9650 9595
rect 9525 9501 9650 9539
rect 10165 9835 10203 9887
rect 10255 9835 10294 9887
rect 8393 9393 8732 9434
rect 8393 9341 8430 9393
rect 8482 9341 8642 9393
rect 8694 9341 8732 9393
rect 8393 9301 8732 9341
rect 8498 5689 8627 9301
rect 7984 5555 8627 5689
rect 7984 4077 8113 5555
rect 8212 3581 8341 4659
rect 9389 3984 9518 4659
rect 9389 3932 9428 3984
rect 9480 3932 9518 3984
rect 9389 3891 9518 3932
rect 8212 3529 8251 3581
rect 8303 3529 8341 3581
rect 8212 3488 8341 3529
rect 9903 3379 10032 4659
rect 10165 4553 10294 9835
rect 11080 3782 11209 4659
rect 11080 3730 11119 3782
rect 11171 3730 11209 3782
rect 11080 3689 11209 3730
rect 9903 3327 9942 3379
rect 9994 3327 10032 3379
rect 9903 3286 10032 3327
rect 11594 3177 11723 4428
rect 11594 3125 11633 3177
rect 11685 3125 11723 3177
rect 11594 3084 11723 3125
rect 8267 212 8396 346
rect 9958 212 10087 346
rect 11649 212 11778 346
<< via2 >>
rect 7346 10820 7402 10822
rect 7346 10768 7348 10820
rect 7348 10768 7400 10820
rect 7400 10768 7402 10820
rect 7346 10766 7402 10768
rect 7346 10602 7402 10604
rect 7346 10550 7348 10602
rect 7348 10550 7400 10602
rect 7400 10550 7402 10602
rect 7346 10548 7402 10550
rect 7346 10384 7402 10386
rect 7346 10332 7348 10384
rect 7348 10332 7400 10384
rect 7400 10332 7402 10384
rect 7346 10330 7402 10332
rect 7785 10820 7841 10822
rect 7785 10768 7787 10820
rect 7787 10768 7839 10820
rect 7839 10768 7841 10820
rect 7785 10766 7841 10768
rect 9169 10763 9225 10765
rect 9169 10711 9171 10763
rect 9171 10711 9223 10763
rect 9223 10711 9225 10763
rect 9169 10709 9225 10711
rect 7785 10602 7841 10604
rect 7785 10550 7787 10602
rect 7787 10550 7839 10602
rect 7839 10550 7841 10602
rect 7785 10548 7841 10550
rect 7785 10384 7841 10386
rect 7785 10332 7787 10384
rect 7787 10332 7839 10384
rect 7839 10332 7841 10384
rect 7785 10330 7841 10332
rect 9169 10545 9225 10547
rect 9169 10493 9171 10545
rect 9171 10493 9223 10545
rect 9223 10493 9225 10545
rect 9169 10491 9225 10493
rect 9169 10327 9225 10329
rect 9169 10275 9171 10327
rect 9171 10275 9223 10327
rect 9223 10275 9225 10327
rect 9169 10273 9225 10275
rect 7346 9797 7402 9799
rect 7346 9745 7348 9797
rect 7348 9745 7400 9797
rect 7400 9745 7402 9797
rect 7346 9743 7402 9745
rect 7346 9579 7402 9581
rect 7346 9527 7348 9579
rect 7348 9527 7400 9579
rect 7400 9527 7402 9579
rect 7346 9525 7402 9527
rect 8532 9856 8588 9858
rect 8532 9804 8534 9856
rect 8534 9804 8586 9856
rect 8586 9804 8588 9856
rect 8532 9802 8588 9804
rect 8532 9638 8588 9640
rect 8532 9586 8534 9638
rect 8534 9586 8586 9638
rect 8586 9586 8588 9638
rect 8532 9584 8588 9586
rect 9560 9811 9616 9813
rect 9560 9759 9562 9811
rect 9562 9759 9614 9811
rect 9614 9759 9616 9811
rect 9560 9757 9616 9759
rect 9560 9593 9616 9595
rect 9560 9541 9562 9593
rect 9562 9541 9614 9593
rect 9614 9541 9616 9593
rect 9560 9539 9616 9541
<< metal3 >>
rect 6791 10822 12165 10971
rect 6791 10766 7346 10822
rect 7402 10766 7785 10822
rect 7841 10766 12165 10822
rect 6791 10765 12165 10766
rect 6791 10709 9169 10765
rect 9225 10709 12165 10765
rect 6791 10604 12165 10709
rect 6791 10548 7346 10604
rect 7402 10548 7785 10604
rect 7841 10548 12165 10604
rect 6791 10547 12165 10548
rect 6791 10491 9169 10547
rect 9225 10491 12165 10547
rect 6791 10386 12165 10491
rect 6791 10330 7346 10386
rect 7402 10330 7785 10386
rect 7841 10330 12165 10386
rect 6791 10329 12165 10330
rect 6791 10273 9169 10329
rect 9225 10273 12165 10329
rect 6791 10019 12165 10273
rect -1 9858 12165 9907
rect -1 9802 8532 9858
rect 8588 9813 12165 9858
rect 8588 9802 9560 9813
rect -1 9799 9560 9802
rect -1 9743 7346 9799
rect 7402 9757 9560 9799
rect 9616 9757 12165 9813
rect 7402 9743 12165 9757
rect -1 9640 12165 9743
rect -1 9584 8532 9640
rect 8588 9595 12165 9640
rect 8588 9584 9560 9595
rect -1 9581 9560 9584
rect -1 9525 7346 9581
rect 7402 9539 9560 9581
rect 9616 9539 12165 9595
rect 7402 9525 12165 9539
rect -1 9194 12165 9525
rect -1 8151 12215 9060
rect -1 5090 12233 7813
rect -1 2234 11985 2916
rect -1 1078 11985 1986
rect 11750 523 11879 656
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_0
timestamp 1666464484
transform 1 0 4563 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_1
timestamp 1666464484
transform 1 0 3891 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_2
timestamp 1666464484
transform 1 0 400 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_3
timestamp 1666464484
transform 1 0 1520 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_4
timestamp 1666464484
transform 1 0 5749 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_5
timestamp 1666464484
transform 1 0 5973 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_6
timestamp 1666464484
transform 1 0 1072 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_7
timestamp 1666464484
transform 1 0 848 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_8
timestamp 1666464484
transform 1 0 4787 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_9
timestamp 1666464484
transform 1 0 3667 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_10
timestamp 1666464484
transform 1 0 5525 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_11
timestamp 1666464484
transform 1 0 6197 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_12
timestamp 1666464484
transform 1 0 2929 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_13
timestamp 1666464484
transform 1 0 2257 0 1 3353
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_14
timestamp 1666464484
transform 1 0 2705 0 1 3151
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_15
timestamp 1666464484
transform 1 0 2481 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_16
timestamp 1666464484
transform 1 0 6421 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_17
timestamp 1666464484
transform 1 0 3153 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_18
timestamp 1666464484
transform 1 0 2033 0 1 4160
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_19
timestamp 1666464484
transform 1 0 5301 0 1 3555
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_20
timestamp 1666464484
transform 1 0 1296 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_21
timestamp 1666464484
transform 1 0 624 0 1 3960
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_22
timestamp 1666464484
transform 1 0 4115 0 1 3756
box 0 0 1 1
use M1_POLY2$$44753964_64x8m81  M1_POLY2$$44753964_64x8m81_23
timestamp 1666464484
transform 1 0 4339 0 1 3151
box 0 0 1 1
use M1_POLY2$$44754988_R270_64x8m81  M1_POLY2$$44754988_R270_64x8m81_0
timestamp 1666464484
transform 0 -1 7324 -1 0 10090
box 0 0 1 1
use M1_POLY24310589983234_64x8m81  M1_POLY24310589983234_64x8m81_0
timestamp 1666464484
transform 1 0 9070 0 1 9417
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1666464484
transform 1 0 8267 0 1 10062
box 0 0 1 1
use M1_POLY24310589983242_64x8m81  M1_POLY24310589983242_64x8m81_0
timestamp 1666464484
transform 1 0 8007 0 1 10386
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_0
timestamp 1666464484
transform -1 0 7291 0 1 10088
box 0 0 1 1
use M2_M1$$34864172_64x8m81  M2_M1$$34864172_64x8m81_1
timestamp 1666464484
transform 1 0 8562 0 1 9367
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1666464484
transform 1 0 8033 0 1 10469
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1666464484
transform 1 0 10229 0 1 9970
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_2
timestamp 1666464484
transform 1 0 8560 0 1 9721
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_3
timestamp 1666464484
transform 1 0 9588 0 1 9676
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_4
timestamp 1666464484
transform 1 0 7374 0 1 9662
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_0
timestamp 1666464484
transform 1 0 9197 0 1 10519
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_1
timestamp 1666464484
transform 1 0 7813 0 1 10576
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_2
timestamp 1666464484
transform 1 0 7374 0 1 10576
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_0
timestamp 1666464484
transform -1 0 11659 0 1 3151
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_1
timestamp 1666464484
transform -1 0 11145 0 1 3756
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_2
timestamp 1666464484
transform -1 0 8277 0 1 3555
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_3
timestamp 1666464484
transform -1 0 9968 0 1 3353
box 0 0 1 1
use M2_M1$$46894124_64x8m81  M2_M1$$46894124_64x8m81_4
timestamp 1666464484
transform -1 0 9454 0 1 3958
box 0 0 1 1
use M2_M1431058998320_64x8m81  M2_M1431058998320_64x8m81_0
timestamp 1666464484
transform 1 0 8211 0 1 10066
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_0
timestamp 1666464484
transform 1 0 8560 0 1 9721
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_1
timestamp 1666464484
transform 1 0 9588 0 1 9676
box 0 0 1 1
use M3_M2$$43368492_64x8m81_0  M3_M2$$43368492_64x8m81_0_2
timestamp 1666464484
transform 1 0 7374 0 1 9662
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_0
timestamp 1666464484
transform 1 0 9197 0 1 10519
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_1
timestamp 1666464484
transform 1 0 7813 0 1 10576
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_2
timestamp 1666464484
transform 1 0 7374 0 1 10576
box 0 0 1 1
use nmos_1p2$$47342636_64x8m81  nmos_1p2$$47342636_64x8m81_0
timestamp 1666464484
transform 1 0 9059 0 1 10236
box -119 -73 177 316
use nmos_5p04310589983260_64x8m81  nmos_5p04310589983260_64x8m81_0
timestamp 1666464484
transform 1 0 7657 0 1 10240
box -88 -44 208 426
use nmos_5p04310589983260_64x8m81  nmos_5p04310589983260_64x8m81_1
timestamp 1666464484
transform 1 0 7433 0 1 10240
box -88 -44 208 426
use pmos_1p2$$47109164_64x8m81  pmos_1p2$$47109164_64x8m81_0
timestamp 1666464484
transform 1 0 8940 0 1 9519
box -239 -120 521 462
use xpredec1_bot_64x8m81  xpredec1_bot_64x8m81_0
timestamp 1666464484
transform 1 0 10222 0 1 632
box -106 -633 1824 8602
use xpredec1_bot_64x8m81  xpredec1_bot_64x8m81_1
timestamp 1666464484
transform 1 0 6841 0 1 632
box -106 -633 1824 8602
use xpredec1_bot_64x8m81  xpredec1_bot_64x8m81_2
timestamp 1666464484
transform 1 0 8531 0 1 632
box -106 -633 1824 8602
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_0
timestamp 1666464484
transform -1 0 4372 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_1
timestamp 1666464484
transform -1 0 6006 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_2
timestamp 1666464484
transform -1 0 2739 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_3
timestamp 1666464484
transform -1 0 1105 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_4
timestamp 1666464484
transform 1 0 4082 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_5
timestamp 1666464484
transform 1 0 5716 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_6
timestamp 1666464484
transform 1 0 2449 0 1 10644
box -144 -10645 1106 327
use xpredec1_xa_64x8m81  xpredec1_xa_64x8m81_7
timestamp 1666464484
transform 1 0 815 0 1 10644
box -144 -10645 1106 327
<< labels >>
rlabel metal3 s 11999 9542 11999 9542 4 vdd
port 1 nsew
rlabel metal3 s 11999 8560 11999 8560 4 vss
port 2 nsew
rlabel metal3 s 11999 6450 11999 6450 4 vdd
port 1 nsew
rlabel metal3 s 11782 1596 11782 1596 4 vdd
port 1 nsew
rlabel metal3 s 11814 2575 11814 2575 4 vss
port 2 nsew
rlabel metal3 s 11814 589 11814 589 4 vss
port 2 nsew
rlabel metal3 s 11999 10557 11999 10557 4 vss
port 2 nsew
rlabel metal2 s 8332 279 8332 279 4 A[2]
port 3 nsew
rlabel metal2 s 7185 10093 7185 10093 4 men
port 4 nsew
rlabel metal2 s 784 10904 784 10904 4 x[7]
port 5 nsew
rlabel metal2 s 1138 10904 1138 10904 4 x[6]
port 6 nsew
rlabel metal2 s 2418 10904 2418 10904 4 x[5]
port 7 nsew
rlabel metal2 s 2780 10904 2780 10904 4 x[4]
port 8 nsew
rlabel metal2 s 4049 10904 4049 10904 4 x[3]
port 9 nsew
rlabel metal2 s 4403 10904 4403 10904 4 x[2]
port 10 nsew
rlabel metal2 s 5710 10904 5710 10904 4 x[1]
port 11 nsew
rlabel metal2 s 6032 10904 6032 10904 4 x[0]
port 12 nsew
rlabel metal2 s 10023 279 10023 279 4 A[1]
port 13 nsew
rlabel metal2 s 11713 279 11713 279 4 A[0]
port 14 nsew
rlabel metal2 s 8033 10573 8033 10573 4 clk
port 15 nsew
<< properties >>
string GDS_END 1097406
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1087726
<< end >>
