magic
tech gf180mcuC
timestamp 1666464484
<< properties >>
string GDS_END 961746
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 961454
<< end >>
