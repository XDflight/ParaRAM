magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 2344 1064
<< mvpmos >>
rect 0 0 120 944
rect 224 0 344 944
rect 448 0 568 944
rect 672 0 792 944
rect 896 0 1016 944
rect 1120 0 1240 944
rect 1344 0 1464 944
rect 1568 0 1688 944
rect 1792 0 1912 944
rect 2016 0 2136 944
<< mvpdiff >>
rect -88 931 0 944
rect -88 885 -75 931
rect -29 885 0 931
rect -88 822 0 885
rect -88 776 -75 822
rect -29 776 0 822
rect -88 713 0 776
rect -88 667 -75 713
rect -29 667 0 713
rect -88 604 0 667
rect -88 558 -75 604
rect -29 558 0 604
rect -88 495 0 558
rect -88 449 -75 495
rect -29 449 0 495
rect -88 386 0 449
rect -88 340 -75 386
rect -29 340 0 386
rect -88 277 0 340
rect -88 231 -75 277
rect -29 231 0 277
rect -88 168 0 231
rect -88 122 -75 168
rect -29 122 0 168
rect -88 59 0 122
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 931 224 944
rect 120 885 149 931
rect 195 885 224 931
rect 120 822 224 885
rect 120 776 149 822
rect 195 776 224 822
rect 120 713 224 776
rect 120 667 149 713
rect 195 667 224 713
rect 120 604 224 667
rect 120 558 149 604
rect 195 558 224 604
rect 120 495 224 558
rect 120 449 149 495
rect 195 449 224 495
rect 120 386 224 449
rect 120 340 149 386
rect 195 340 224 386
rect 120 277 224 340
rect 120 231 149 277
rect 195 231 224 277
rect 120 168 224 231
rect 120 122 149 168
rect 195 122 224 168
rect 120 59 224 122
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 931 448 944
rect 344 885 373 931
rect 419 885 448 931
rect 344 822 448 885
rect 344 776 373 822
rect 419 776 448 822
rect 344 713 448 776
rect 344 667 373 713
rect 419 667 448 713
rect 344 604 448 667
rect 344 558 373 604
rect 419 558 448 604
rect 344 495 448 558
rect 344 449 373 495
rect 419 449 448 495
rect 344 386 448 449
rect 344 340 373 386
rect 419 340 448 386
rect 344 277 448 340
rect 344 231 373 277
rect 419 231 448 277
rect 344 168 448 231
rect 344 122 373 168
rect 419 122 448 168
rect 344 59 448 122
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 931 672 944
rect 568 885 597 931
rect 643 885 672 931
rect 568 822 672 885
rect 568 776 597 822
rect 643 776 672 822
rect 568 713 672 776
rect 568 667 597 713
rect 643 667 672 713
rect 568 604 672 667
rect 568 558 597 604
rect 643 558 672 604
rect 568 495 672 558
rect 568 449 597 495
rect 643 449 672 495
rect 568 386 672 449
rect 568 340 597 386
rect 643 340 672 386
rect 568 277 672 340
rect 568 231 597 277
rect 643 231 672 277
rect 568 168 672 231
rect 568 122 597 168
rect 643 122 672 168
rect 568 59 672 122
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 931 896 944
rect 792 885 821 931
rect 867 885 896 931
rect 792 822 896 885
rect 792 776 821 822
rect 867 776 896 822
rect 792 713 896 776
rect 792 667 821 713
rect 867 667 896 713
rect 792 604 896 667
rect 792 558 821 604
rect 867 558 896 604
rect 792 495 896 558
rect 792 449 821 495
rect 867 449 896 495
rect 792 386 896 449
rect 792 340 821 386
rect 867 340 896 386
rect 792 277 896 340
rect 792 231 821 277
rect 867 231 896 277
rect 792 168 896 231
rect 792 122 821 168
rect 867 122 896 168
rect 792 59 896 122
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 931 1120 944
rect 1016 885 1045 931
rect 1091 885 1120 931
rect 1016 822 1120 885
rect 1016 776 1045 822
rect 1091 776 1120 822
rect 1016 713 1120 776
rect 1016 667 1045 713
rect 1091 667 1120 713
rect 1016 604 1120 667
rect 1016 558 1045 604
rect 1091 558 1120 604
rect 1016 495 1120 558
rect 1016 449 1045 495
rect 1091 449 1120 495
rect 1016 386 1120 449
rect 1016 340 1045 386
rect 1091 340 1120 386
rect 1016 277 1120 340
rect 1016 231 1045 277
rect 1091 231 1120 277
rect 1016 168 1120 231
rect 1016 122 1045 168
rect 1091 122 1120 168
rect 1016 59 1120 122
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 931 1344 944
rect 1240 885 1269 931
rect 1315 885 1344 931
rect 1240 822 1344 885
rect 1240 776 1269 822
rect 1315 776 1344 822
rect 1240 713 1344 776
rect 1240 667 1269 713
rect 1315 667 1344 713
rect 1240 604 1344 667
rect 1240 558 1269 604
rect 1315 558 1344 604
rect 1240 495 1344 558
rect 1240 449 1269 495
rect 1315 449 1344 495
rect 1240 386 1344 449
rect 1240 340 1269 386
rect 1315 340 1344 386
rect 1240 277 1344 340
rect 1240 231 1269 277
rect 1315 231 1344 277
rect 1240 168 1344 231
rect 1240 122 1269 168
rect 1315 122 1344 168
rect 1240 59 1344 122
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 931 1568 944
rect 1464 885 1493 931
rect 1539 885 1568 931
rect 1464 822 1568 885
rect 1464 776 1493 822
rect 1539 776 1568 822
rect 1464 713 1568 776
rect 1464 667 1493 713
rect 1539 667 1568 713
rect 1464 604 1568 667
rect 1464 558 1493 604
rect 1539 558 1568 604
rect 1464 495 1568 558
rect 1464 449 1493 495
rect 1539 449 1568 495
rect 1464 386 1568 449
rect 1464 340 1493 386
rect 1539 340 1568 386
rect 1464 277 1568 340
rect 1464 231 1493 277
rect 1539 231 1568 277
rect 1464 168 1568 231
rect 1464 122 1493 168
rect 1539 122 1568 168
rect 1464 59 1568 122
rect 1464 13 1493 59
rect 1539 13 1568 59
rect 1464 0 1568 13
rect 1688 931 1792 944
rect 1688 885 1717 931
rect 1763 885 1792 931
rect 1688 822 1792 885
rect 1688 776 1717 822
rect 1763 776 1792 822
rect 1688 713 1792 776
rect 1688 667 1717 713
rect 1763 667 1792 713
rect 1688 604 1792 667
rect 1688 558 1717 604
rect 1763 558 1792 604
rect 1688 495 1792 558
rect 1688 449 1717 495
rect 1763 449 1792 495
rect 1688 386 1792 449
rect 1688 340 1717 386
rect 1763 340 1792 386
rect 1688 277 1792 340
rect 1688 231 1717 277
rect 1763 231 1792 277
rect 1688 168 1792 231
rect 1688 122 1717 168
rect 1763 122 1792 168
rect 1688 59 1792 122
rect 1688 13 1717 59
rect 1763 13 1792 59
rect 1688 0 1792 13
rect 1912 931 2016 944
rect 1912 885 1941 931
rect 1987 885 2016 931
rect 1912 822 2016 885
rect 1912 776 1941 822
rect 1987 776 2016 822
rect 1912 713 2016 776
rect 1912 667 1941 713
rect 1987 667 2016 713
rect 1912 604 2016 667
rect 1912 558 1941 604
rect 1987 558 2016 604
rect 1912 495 2016 558
rect 1912 449 1941 495
rect 1987 449 2016 495
rect 1912 386 2016 449
rect 1912 340 1941 386
rect 1987 340 2016 386
rect 1912 277 2016 340
rect 1912 231 1941 277
rect 1987 231 2016 277
rect 1912 168 2016 231
rect 1912 122 1941 168
rect 1987 122 2016 168
rect 1912 59 2016 122
rect 1912 13 1941 59
rect 1987 13 2016 59
rect 1912 0 2016 13
rect 2136 931 2224 944
rect 2136 885 2165 931
rect 2211 885 2224 931
rect 2136 822 2224 885
rect 2136 776 2165 822
rect 2211 776 2224 822
rect 2136 713 2224 776
rect 2136 667 2165 713
rect 2211 667 2224 713
rect 2136 604 2224 667
rect 2136 558 2165 604
rect 2211 558 2224 604
rect 2136 495 2224 558
rect 2136 449 2165 495
rect 2211 449 2224 495
rect 2136 386 2224 449
rect 2136 340 2165 386
rect 2211 340 2224 386
rect 2136 277 2224 340
rect 2136 231 2165 277
rect 2211 231 2224 277
rect 2136 168 2224 231
rect 2136 122 2165 168
rect 2211 122 2224 168
rect 2136 59 2224 122
rect 2136 13 2165 59
rect 2211 13 2224 59
rect 2136 0 2224 13
<< mvpdiffc >>
rect -75 885 -29 931
rect -75 776 -29 822
rect -75 667 -29 713
rect -75 558 -29 604
rect -75 449 -29 495
rect -75 340 -29 386
rect -75 231 -29 277
rect -75 122 -29 168
rect -75 13 -29 59
rect 149 885 195 931
rect 149 776 195 822
rect 149 667 195 713
rect 149 558 195 604
rect 149 449 195 495
rect 149 340 195 386
rect 149 231 195 277
rect 149 122 195 168
rect 149 13 195 59
rect 373 885 419 931
rect 373 776 419 822
rect 373 667 419 713
rect 373 558 419 604
rect 373 449 419 495
rect 373 340 419 386
rect 373 231 419 277
rect 373 122 419 168
rect 373 13 419 59
rect 597 885 643 931
rect 597 776 643 822
rect 597 667 643 713
rect 597 558 643 604
rect 597 449 643 495
rect 597 340 643 386
rect 597 231 643 277
rect 597 122 643 168
rect 597 13 643 59
rect 821 885 867 931
rect 821 776 867 822
rect 821 667 867 713
rect 821 558 867 604
rect 821 449 867 495
rect 821 340 867 386
rect 821 231 867 277
rect 821 122 867 168
rect 821 13 867 59
rect 1045 885 1091 931
rect 1045 776 1091 822
rect 1045 667 1091 713
rect 1045 558 1091 604
rect 1045 449 1091 495
rect 1045 340 1091 386
rect 1045 231 1091 277
rect 1045 122 1091 168
rect 1045 13 1091 59
rect 1269 885 1315 931
rect 1269 776 1315 822
rect 1269 667 1315 713
rect 1269 558 1315 604
rect 1269 449 1315 495
rect 1269 340 1315 386
rect 1269 231 1315 277
rect 1269 122 1315 168
rect 1269 13 1315 59
rect 1493 885 1539 931
rect 1493 776 1539 822
rect 1493 667 1539 713
rect 1493 558 1539 604
rect 1493 449 1539 495
rect 1493 340 1539 386
rect 1493 231 1539 277
rect 1493 122 1539 168
rect 1493 13 1539 59
rect 1717 885 1763 931
rect 1717 776 1763 822
rect 1717 667 1763 713
rect 1717 558 1763 604
rect 1717 449 1763 495
rect 1717 340 1763 386
rect 1717 231 1763 277
rect 1717 122 1763 168
rect 1717 13 1763 59
rect 1941 885 1987 931
rect 1941 776 1987 822
rect 1941 667 1987 713
rect 1941 558 1987 604
rect 1941 449 1987 495
rect 1941 340 1987 386
rect 1941 231 1987 277
rect 1941 122 1987 168
rect 1941 13 1987 59
rect 2165 885 2211 931
rect 2165 776 2211 822
rect 2165 667 2211 713
rect 2165 558 2211 604
rect 2165 449 2211 495
rect 2165 340 2211 386
rect 2165 231 2211 277
rect 2165 122 2211 168
rect 2165 13 2211 59
<< polysilicon >>
rect 0 944 120 988
rect 224 944 344 988
rect 448 944 568 988
rect 672 944 792 988
rect 896 944 1016 988
rect 1120 944 1240 988
rect 1344 944 1464 988
rect 1568 944 1688 988
rect 1792 944 1912 988
rect 2016 944 2136 988
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
<< metal1 >>
rect -75 931 -29 944
rect -75 822 -29 885
rect -75 713 -29 776
rect -75 604 -29 667
rect -75 495 -29 558
rect -75 386 -29 449
rect -75 277 -29 340
rect -75 168 -29 231
rect -75 59 -29 122
rect -75 0 -29 13
rect 149 931 195 944
rect 149 822 195 885
rect 149 713 195 776
rect 149 604 195 667
rect 149 495 195 558
rect 149 386 195 449
rect 149 277 195 340
rect 149 168 195 231
rect 149 59 195 122
rect 149 0 195 13
rect 373 931 419 944
rect 373 822 419 885
rect 373 713 419 776
rect 373 604 419 667
rect 373 495 419 558
rect 373 386 419 449
rect 373 277 419 340
rect 373 168 419 231
rect 373 59 419 122
rect 373 0 419 13
rect 597 931 643 944
rect 597 822 643 885
rect 597 713 643 776
rect 597 604 643 667
rect 597 495 643 558
rect 597 386 643 449
rect 597 277 643 340
rect 597 168 643 231
rect 597 59 643 122
rect 597 0 643 13
rect 821 931 867 944
rect 821 822 867 885
rect 821 713 867 776
rect 821 604 867 667
rect 821 495 867 558
rect 821 386 867 449
rect 821 277 867 340
rect 821 168 867 231
rect 821 59 867 122
rect 821 0 867 13
rect 1045 931 1091 944
rect 1045 822 1091 885
rect 1045 713 1091 776
rect 1045 604 1091 667
rect 1045 495 1091 558
rect 1045 386 1091 449
rect 1045 277 1091 340
rect 1045 168 1091 231
rect 1045 59 1091 122
rect 1045 0 1091 13
rect 1269 931 1315 944
rect 1269 822 1315 885
rect 1269 713 1315 776
rect 1269 604 1315 667
rect 1269 495 1315 558
rect 1269 386 1315 449
rect 1269 277 1315 340
rect 1269 168 1315 231
rect 1269 59 1315 122
rect 1269 0 1315 13
rect 1493 931 1539 944
rect 1493 822 1539 885
rect 1493 713 1539 776
rect 1493 604 1539 667
rect 1493 495 1539 558
rect 1493 386 1539 449
rect 1493 277 1539 340
rect 1493 168 1539 231
rect 1493 59 1539 122
rect 1493 0 1539 13
rect 1717 931 1763 944
rect 1717 822 1763 885
rect 1717 713 1763 776
rect 1717 604 1763 667
rect 1717 495 1763 558
rect 1717 386 1763 449
rect 1717 277 1763 340
rect 1717 168 1763 231
rect 1717 59 1763 122
rect 1717 0 1763 13
rect 1941 931 1987 944
rect 1941 822 1987 885
rect 1941 713 1987 776
rect 1941 604 1987 667
rect 1941 495 1987 558
rect 1941 386 1987 449
rect 1941 277 1987 340
rect 1941 168 1987 231
rect 1941 59 1987 122
rect 1941 0 1987 13
rect 2165 931 2211 944
rect 2165 822 2211 885
rect 2165 713 2211 776
rect 2165 604 2211 667
rect 2165 495 2211 558
rect 2165 386 2211 449
rect 2165 277 2211 340
rect 2165 168 2211 231
rect 2165 59 2211 122
rect 2165 0 2211 13
<< labels >>
flabel metal1 s -52 472 -52 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 2188 472 2188 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 472 172 472 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 472 396 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 472 620 472 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 472 844 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 472 1068 472 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 472 1292 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 472 1516 472 0 FreeSans 400 0 0 0 D
flabel metal1 s 1740 472 1740 472 0 FreeSans 400 0 0 0 S
flabel metal1 s 1964 472 1964 472 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 322598
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 311864
<< end >>
