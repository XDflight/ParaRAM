magic
tech gf180mcuC
magscale 1 5
timestamp 1667635171
<< obsm1 >>
rect 672 855 89320 58561
<< metal2 >>
rect 672 59600 728 60000
rect 1456 59600 1512 60000
rect 2240 59600 2296 60000
rect 3024 59600 3080 60000
rect 3808 59600 3864 60000
rect 4592 59600 4648 60000
rect 5376 59600 5432 60000
rect 6160 59600 6216 60000
rect 6944 59600 7000 60000
rect 7728 59600 7784 60000
rect 8512 59600 8568 60000
rect 9296 59600 9352 60000
rect 10080 59600 10136 60000
rect 10864 59600 10920 60000
rect 11648 59600 11704 60000
rect 12432 59600 12488 60000
rect 13216 59600 13272 60000
rect 14000 59600 14056 60000
rect 14784 59600 14840 60000
rect 15568 59600 15624 60000
rect 16352 59600 16408 60000
rect 17136 59600 17192 60000
rect 17920 59600 17976 60000
rect 18704 59600 18760 60000
rect 19488 59600 19544 60000
rect 20272 59600 20328 60000
rect 21056 59600 21112 60000
rect 21840 59600 21896 60000
rect 22624 59600 22680 60000
rect 23408 59600 23464 60000
rect 24192 59600 24248 60000
rect 24976 59600 25032 60000
rect 25760 59600 25816 60000
rect 26544 59600 26600 60000
rect 27328 59600 27384 60000
rect 28112 59600 28168 60000
rect 28896 59600 28952 60000
rect 29680 59600 29736 60000
rect 30464 59600 30520 60000
rect 31248 59600 31304 60000
rect 32032 59600 32088 60000
rect 32816 59600 32872 60000
rect 33600 59600 33656 60000
rect 34384 59600 34440 60000
rect 35168 59600 35224 60000
rect 35952 59600 36008 60000
rect 36736 59600 36792 60000
rect 37520 59600 37576 60000
rect 38304 59600 38360 60000
rect 39088 59600 39144 60000
rect 39872 59600 39928 60000
rect 40656 59600 40712 60000
rect 41440 59600 41496 60000
rect 42224 59600 42280 60000
rect 43008 59600 43064 60000
rect 43792 59600 43848 60000
rect 44576 59600 44632 60000
rect 45360 59600 45416 60000
rect 46144 59600 46200 60000
rect 46928 59600 46984 60000
rect 47712 59600 47768 60000
rect 48496 59600 48552 60000
rect 49280 59600 49336 60000
rect 50064 59600 50120 60000
rect 50848 59600 50904 60000
rect 51632 59600 51688 60000
rect 52416 59600 52472 60000
rect 53200 59600 53256 60000
rect 53984 59600 54040 60000
rect 54768 59600 54824 60000
rect 55552 59600 55608 60000
rect 56336 59600 56392 60000
rect 57120 59600 57176 60000
rect 57904 59600 57960 60000
rect 58688 59600 58744 60000
rect 59472 59600 59528 60000
rect 60256 59600 60312 60000
rect 61040 59600 61096 60000
rect 61824 59600 61880 60000
rect 62608 59600 62664 60000
rect 63392 59600 63448 60000
rect 64176 59600 64232 60000
rect 64960 59600 65016 60000
rect 65744 59600 65800 60000
rect 66528 59600 66584 60000
rect 67312 59600 67368 60000
rect 68096 59600 68152 60000
rect 68880 59600 68936 60000
rect 69664 59600 69720 60000
rect 70448 59600 70504 60000
rect 71232 59600 71288 60000
rect 72016 59600 72072 60000
rect 72800 59600 72856 60000
rect 73584 59600 73640 60000
rect 74368 59600 74424 60000
rect 75152 59600 75208 60000
rect 75936 59600 75992 60000
rect 76720 59600 76776 60000
rect 77504 59600 77560 60000
rect 78288 59600 78344 60000
rect 79072 59600 79128 60000
rect 79856 59600 79912 60000
rect 80640 59600 80696 60000
rect 81424 59600 81480 60000
rect 82208 59600 82264 60000
rect 82992 59600 83048 60000
rect 83776 59600 83832 60000
rect 84560 59600 84616 60000
rect 85344 59600 85400 60000
rect 86128 59600 86184 60000
rect 86912 59600 86968 60000
rect 87696 59600 87752 60000
rect 88480 59600 88536 60000
rect 89264 59600 89320 60000
rect 3640 0 3696 400
rect 3808 0 3864 400
rect 3976 0 4032 400
rect 4144 0 4200 400
rect 4312 0 4368 400
rect 4480 0 4536 400
rect 4648 0 4704 400
rect 4816 0 4872 400
rect 4984 0 5040 400
rect 5152 0 5208 400
rect 5320 0 5376 400
rect 5488 0 5544 400
rect 5656 0 5712 400
rect 5824 0 5880 400
rect 5992 0 6048 400
rect 6160 0 6216 400
rect 6328 0 6384 400
rect 6496 0 6552 400
rect 6664 0 6720 400
rect 6832 0 6888 400
rect 7000 0 7056 400
rect 7168 0 7224 400
rect 7336 0 7392 400
rect 7504 0 7560 400
rect 7672 0 7728 400
rect 7840 0 7896 400
rect 8008 0 8064 400
rect 8176 0 8232 400
rect 8344 0 8400 400
rect 8512 0 8568 400
rect 8680 0 8736 400
rect 8848 0 8904 400
rect 9016 0 9072 400
rect 9184 0 9240 400
rect 9352 0 9408 400
rect 9520 0 9576 400
rect 9688 0 9744 400
rect 9856 0 9912 400
rect 10024 0 10080 400
rect 10192 0 10248 400
rect 10360 0 10416 400
rect 10528 0 10584 400
rect 10696 0 10752 400
rect 10864 0 10920 400
rect 11032 0 11088 400
rect 11200 0 11256 400
rect 11368 0 11424 400
rect 11536 0 11592 400
rect 11704 0 11760 400
rect 11872 0 11928 400
rect 12040 0 12096 400
rect 12208 0 12264 400
rect 12376 0 12432 400
rect 12544 0 12600 400
rect 12712 0 12768 400
rect 12880 0 12936 400
rect 13048 0 13104 400
rect 13216 0 13272 400
rect 13384 0 13440 400
rect 13552 0 13608 400
rect 13720 0 13776 400
rect 13888 0 13944 400
rect 14056 0 14112 400
rect 14224 0 14280 400
rect 14392 0 14448 400
rect 14560 0 14616 400
rect 14728 0 14784 400
rect 14896 0 14952 400
rect 15064 0 15120 400
rect 15232 0 15288 400
rect 15400 0 15456 400
rect 15568 0 15624 400
rect 15736 0 15792 400
rect 15904 0 15960 400
rect 16072 0 16128 400
rect 16240 0 16296 400
rect 16408 0 16464 400
rect 16576 0 16632 400
rect 16744 0 16800 400
rect 16912 0 16968 400
rect 17080 0 17136 400
rect 17248 0 17304 400
rect 17416 0 17472 400
rect 17584 0 17640 400
rect 17752 0 17808 400
rect 17920 0 17976 400
rect 18088 0 18144 400
rect 18256 0 18312 400
rect 18424 0 18480 400
rect 18592 0 18648 400
rect 18760 0 18816 400
rect 18928 0 18984 400
rect 19096 0 19152 400
rect 19264 0 19320 400
rect 19432 0 19488 400
rect 19600 0 19656 400
rect 19768 0 19824 400
rect 19936 0 19992 400
rect 20104 0 20160 400
rect 20272 0 20328 400
rect 20440 0 20496 400
rect 20608 0 20664 400
rect 20776 0 20832 400
rect 20944 0 21000 400
rect 21112 0 21168 400
rect 21280 0 21336 400
rect 21448 0 21504 400
rect 21616 0 21672 400
rect 21784 0 21840 400
rect 21952 0 22008 400
rect 22120 0 22176 400
rect 22288 0 22344 400
rect 22456 0 22512 400
rect 22624 0 22680 400
rect 22792 0 22848 400
rect 22960 0 23016 400
rect 23128 0 23184 400
rect 23296 0 23352 400
rect 23464 0 23520 400
rect 23632 0 23688 400
rect 23800 0 23856 400
rect 23968 0 24024 400
rect 24136 0 24192 400
rect 24304 0 24360 400
rect 24472 0 24528 400
rect 24640 0 24696 400
rect 24808 0 24864 400
rect 24976 0 25032 400
rect 25144 0 25200 400
rect 25312 0 25368 400
rect 25480 0 25536 400
rect 25648 0 25704 400
rect 25816 0 25872 400
rect 25984 0 26040 400
rect 26152 0 26208 400
rect 26320 0 26376 400
rect 26488 0 26544 400
rect 26656 0 26712 400
rect 26824 0 26880 400
rect 26992 0 27048 400
rect 27160 0 27216 400
rect 27328 0 27384 400
rect 27496 0 27552 400
rect 27664 0 27720 400
rect 27832 0 27888 400
rect 28000 0 28056 400
rect 28168 0 28224 400
rect 28336 0 28392 400
rect 28504 0 28560 400
rect 28672 0 28728 400
rect 28840 0 28896 400
rect 29008 0 29064 400
rect 29176 0 29232 400
rect 29344 0 29400 400
rect 29512 0 29568 400
rect 29680 0 29736 400
rect 29848 0 29904 400
rect 30016 0 30072 400
rect 30184 0 30240 400
rect 30352 0 30408 400
rect 30520 0 30576 400
rect 30688 0 30744 400
rect 30856 0 30912 400
rect 31024 0 31080 400
rect 31192 0 31248 400
rect 31360 0 31416 400
rect 31528 0 31584 400
rect 31696 0 31752 400
rect 31864 0 31920 400
rect 32032 0 32088 400
rect 32200 0 32256 400
rect 32368 0 32424 400
rect 32536 0 32592 400
rect 32704 0 32760 400
rect 32872 0 32928 400
rect 33040 0 33096 400
rect 33208 0 33264 400
rect 33376 0 33432 400
rect 33544 0 33600 400
rect 33712 0 33768 400
rect 33880 0 33936 400
rect 34048 0 34104 400
rect 34216 0 34272 400
rect 34384 0 34440 400
rect 34552 0 34608 400
rect 34720 0 34776 400
rect 34888 0 34944 400
rect 35056 0 35112 400
rect 35224 0 35280 400
rect 35392 0 35448 400
rect 35560 0 35616 400
rect 35728 0 35784 400
rect 35896 0 35952 400
rect 36064 0 36120 400
rect 36232 0 36288 400
rect 36400 0 36456 400
rect 36568 0 36624 400
rect 36736 0 36792 400
rect 36904 0 36960 400
rect 37072 0 37128 400
rect 37240 0 37296 400
rect 37408 0 37464 400
rect 37576 0 37632 400
rect 37744 0 37800 400
rect 37912 0 37968 400
rect 38080 0 38136 400
rect 38248 0 38304 400
rect 38416 0 38472 400
rect 38584 0 38640 400
rect 38752 0 38808 400
rect 38920 0 38976 400
rect 39088 0 39144 400
rect 39256 0 39312 400
rect 39424 0 39480 400
rect 39592 0 39648 400
rect 39760 0 39816 400
rect 39928 0 39984 400
rect 40096 0 40152 400
rect 40264 0 40320 400
rect 40432 0 40488 400
rect 40600 0 40656 400
rect 40768 0 40824 400
rect 40936 0 40992 400
rect 41104 0 41160 400
rect 41272 0 41328 400
rect 41440 0 41496 400
rect 41608 0 41664 400
rect 41776 0 41832 400
rect 41944 0 42000 400
rect 42112 0 42168 400
rect 42280 0 42336 400
rect 42448 0 42504 400
rect 42616 0 42672 400
rect 42784 0 42840 400
rect 42952 0 43008 400
rect 43120 0 43176 400
rect 43288 0 43344 400
rect 43456 0 43512 400
rect 43624 0 43680 400
rect 43792 0 43848 400
rect 43960 0 44016 400
rect 44128 0 44184 400
rect 44296 0 44352 400
rect 44464 0 44520 400
rect 44632 0 44688 400
rect 44800 0 44856 400
rect 44968 0 45024 400
rect 45136 0 45192 400
rect 45304 0 45360 400
rect 45472 0 45528 400
rect 45640 0 45696 400
rect 45808 0 45864 400
rect 45976 0 46032 400
rect 46144 0 46200 400
rect 46312 0 46368 400
rect 46480 0 46536 400
rect 46648 0 46704 400
rect 46816 0 46872 400
rect 46984 0 47040 400
rect 47152 0 47208 400
rect 47320 0 47376 400
rect 47488 0 47544 400
rect 47656 0 47712 400
rect 47824 0 47880 400
rect 47992 0 48048 400
rect 48160 0 48216 400
rect 48328 0 48384 400
rect 48496 0 48552 400
rect 48664 0 48720 400
rect 48832 0 48888 400
rect 49000 0 49056 400
rect 49168 0 49224 400
rect 49336 0 49392 400
rect 49504 0 49560 400
rect 49672 0 49728 400
rect 49840 0 49896 400
rect 50008 0 50064 400
rect 50176 0 50232 400
rect 50344 0 50400 400
rect 50512 0 50568 400
rect 50680 0 50736 400
rect 50848 0 50904 400
rect 51016 0 51072 400
rect 51184 0 51240 400
rect 51352 0 51408 400
rect 51520 0 51576 400
rect 51688 0 51744 400
rect 51856 0 51912 400
rect 52024 0 52080 400
rect 52192 0 52248 400
rect 52360 0 52416 400
rect 52528 0 52584 400
rect 52696 0 52752 400
rect 52864 0 52920 400
rect 53032 0 53088 400
rect 53200 0 53256 400
rect 53368 0 53424 400
rect 53536 0 53592 400
rect 53704 0 53760 400
rect 53872 0 53928 400
rect 54040 0 54096 400
rect 54208 0 54264 400
rect 54376 0 54432 400
rect 54544 0 54600 400
rect 54712 0 54768 400
rect 54880 0 54936 400
rect 55048 0 55104 400
rect 55216 0 55272 400
rect 55384 0 55440 400
rect 55552 0 55608 400
rect 55720 0 55776 400
rect 55888 0 55944 400
rect 56056 0 56112 400
rect 56224 0 56280 400
rect 56392 0 56448 400
rect 56560 0 56616 400
rect 56728 0 56784 400
rect 56896 0 56952 400
rect 57064 0 57120 400
rect 57232 0 57288 400
rect 57400 0 57456 400
rect 57568 0 57624 400
rect 57736 0 57792 400
rect 57904 0 57960 400
rect 58072 0 58128 400
rect 58240 0 58296 400
rect 58408 0 58464 400
rect 58576 0 58632 400
rect 58744 0 58800 400
rect 58912 0 58968 400
rect 59080 0 59136 400
rect 59248 0 59304 400
rect 59416 0 59472 400
rect 59584 0 59640 400
rect 59752 0 59808 400
rect 59920 0 59976 400
rect 60088 0 60144 400
rect 60256 0 60312 400
rect 60424 0 60480 400
rect 60592 0 60648 400
rect 60760 0 60816 400
rect 60928 0 60984 400
rect 61096 0 61152 400
rect 61264 0 61320 400
rect 61432 0 61488 400
rect 61600 0 61656 400
rect 61768 0 61824 400
rect 61936 0 61992 400
rect 62104 0 62160 400
rect 62272 0 62328 400
rect 62440 0 62496 400
rect 62608 0 62664 400
rect 62776 0 62832 400
rect 62944 0 63000 400
rect 63112 0 63168 400
rect 63280 0 63336 400
rect 63448 0 63504 400
rect 63616 0 63672 400
rect 63784 0 63840 400
rect 63952 0 64008 400
rect 64120 0 64176 400
rect 64288 0 64344 400
rect 64456 0 64512 400
rect 64624 0 64680 400
rect 64792 0 64848 400
rect 64960 0 65016 400
rect 65128 0 65184 400
rect 65296 0 65352 400
rect 65464 0 65520 400
rect 65632 0 65688 400
rect 65800 0 65856 400
rect 65968 0 66024 400
rect 66136 0 66192 400
rect 66304 0 66360 400
rect 66472 0 66528 400
rect 66640 0 66696 400
rect 66808 0 66864 400
rect 66976 0 67032 400
rect 67144 0 67200 400
rect 67312 0 67368 400
rect 67480 0 67536 400
rect 67648 0 67704 400
rect 67816 0 67872 400
rect 67984 0 68040 400
rect 68152 0 68208 400
rect 68320 0 68376 400
rect 68488 0 68544 400
rect 68656 0 68712 400
rect 68824 0 68880 400
rect 68992 0 69048 400
rect 69160 0 69216 400
rect 69328 0 69384 400
rect 69496 0 69552 400
rect 69664 0 69720 400
rect 69832 0 69888 400
rect 70000 0 70056 400
rect 70168 0 70224 400
rect 70336 0 70392 400
rect 70504 0 70560 400
rect 70672 0 70728 400
rect 70840 0 70896 400
rect 71008 0 71064 400
rect 71176 0 71232 400
rect 71344 0 71400 400
rect 71512 0 71568 400
rect 71680 0 71736 400
rect 71848 0 71904 400
rect 72016 0 72072 400
rect 72184 0 72240 400
rect 72352 0 72408 400
rect 72520 0 72576 400
rect 72688 0 72744 400
rect 72856 0 72912 400
rect 73024 0 73080 400
rect 73192 0 73248 400
rect 73360 0 73416 400
rect 73528 0 73584 400
rect 73696 0 73752 400
rect 73864 0 73920 400
rect 74032 0 74088 400
rect 74200 0 74256 400
rect 74368 0 74424 400
rect 74536 0 74592 400
rect 74704 0 74760 400
rect 74872 0 74928 400
rect 75040 0 75096 400
rect 75208 0 75264 400
rect 75376 0 75432 400
rect 75544 0 75600 400
rect 75712 0 75768 400
rect 75880 0 75936 400
rect 76048 0 76104 400
rect 76216 0 76272 400
rect 76384 0 76440 400
rect 76552 0 76608 400
rect 76720 0 76776 400
rect 76888 0 76944 400
rect 77056 0 77112 400
rect 77224 0 77280 400
rect 77392 0 77448 400
rect 77560 0 77616 400
rect 77728 0 77784 400
rect 77896 0 77952 400
rect 78064 0 78120 400
rect 78232 0 78288 400
rect 78400 0 78456 400
rect 78568 0 78624 400
rect 78736 0 78792 400
rect 78904 0 78960 400
rect 79072 0 79128 400
rect 79240 0 79296 400
rect 79408 0 79464 400
rect 79576 0 79632 400
rect 79744 0 79800 400
rect 79912 0 79968 400
rect 80080 0 80136 400
rect 80248 0 80304 400
rect 80416 0 80472 400
rect 80584 0 80640 400
rect 80752 0 80808 400
rect 80920 0 80976 400
rect 81088 0 81144 400
rect 81256 0 81312 400
rect 81424 0 81480 400
rect 81592 0 81648 400
rect 81760 0 81816 400
rect 81928 0 81984 400
rect 82096 0 82152 400
rect 82264 0 82320 400
rect 82432 0 82488 400
rect 82600 0 82656 400
rect 82768 0 82824 400
rect 82936 0 82992 400
rect 83104 0 83160 400
rect 83272 0 83328 400
rect 83440 0 83496 400
rect 83608 0 83664 400
rect 83776 0 83832 400
rect 83944 0 84000 400
rect 84112 0 84168 400
rect 84280 0 84336 400
rect 84448 0 84504 400
rect 84616 0 84672 400
rect 84784 0 84840 400
rect 84952 0 85008 400
rect 85120 0 85176 400
rect 85288 0 85344 400
rect 85456 0 85512 400
rect 85624 0 85680 400
rect 85792 0 85848 400
rect 85960 0 86016 400
rect 86128 0 86184 400
rect 86296 0 86352 400
<< obsm2 >>
rect 1542 59570 2210 59600
rect 2326 59570 2994 59600
rect 3110 59570 3778 59600
rect 3894 59570 4562 59600
rect 4678 59570 5346 59600
rect 5462 59570 6130 59600
rect 6246 59570 6914 59600
rect 7030 59570 7698 59600
rect 7814 59570 8482 59600
rect 8598 59570 9266 59600
rect 9382 59570 10050 59600
rect 10166 59570 10834 59600
rect 10950 59570 11618 59600
rect 11734 59570 12402 59600
rect 12518 59570 13186 59600
rect 13302 59570 13970 59600
rect 14086 59570 14754 59600
rect 14870 59570 15538 59600
rect 15654 59570 16322 59600
rect 16438 59570 17106 59600
rect 17222 59570 17890 59600
rect 18006 59570 18674 59600
rect 18790 59570 19458 59600
rect 19574 59570 20242 59600
rect 20358 59570 21026 59600
rect 21142 59570 21810 59600
rect 21926 59570 22594 59600
rect 22710 59570 23378 59600
rect 23494 59570 24162 59600
rect 24278 59570 24946 59600
rect 25062 59570 25730 59600
rect 25846 59570 26514 59600
rect 26630 59570 27298 59600
rect 27414 59570 28082 59600
rect 28198 59570 28866 59600
rect 28982 59570 29650 59600
rect 29766 59570 30434 59600
rect 30550 59570 31218 59600
rect 31334 59570 32002 59600
rect 32118 59570 32786 59600
rect 32902 59570 33570 59600
rect 33686 59570 34354 59600
rect 34470 59570 35138 59600
rect 35254 59570 35922 59600
rect 36038 59570 36706 59600
rect 36822 59570 37490 59600
rect 37606 59570 38274 59600
rect 38390 59570 39058 59600
rect 39174 59570 39842 59600
rect 39958 59570 40626 59600
rect 40742 59570 41410 59600
rect 41526 59570 42194 59600
rect 42310 59570 42978 59600
rect 43094 59570 43762 59600
rect 43878 59570 44546 59600
rect 44662 59570 45330 59600
rect 45446 59570 46114 59600
rect 46230 59570 46898 59600
rect 47014 59570 47682 59600
rect 47798 59570 48466 59600
rect 48582 59570 49250 59600
rect 49366 59570 50034 59600
rect 50150 59570 50818 59600
rect 50934 59570 51602 59600
rect 51718 59570 52386 59600
rect 52502 59570 53170 59600
rect 53286 59570 53954 59600
rect 54070 59570 54738 59600
rect 54854 59570 55522 59600
rect 55638 59570 56306 59600
rect 56422 59570 57090 59600
rect 57206 59570 57874 59600
rect 57990 59570 58658 59600
rect 58774 59570 59442 59600
rect 59558 59570 60226 59600
rect 60342 59570 61010 59600
rect 61126 59570 61794 59600
rect 61910 59570 62578 59600
rect 62694 59570 63362 59600
rect 63478 59570 64146 59600
rect 64262 59570 64930 59600
rect 65046 59570 65714 59600
rect 65830 59570 66498 59600
rect 66614 59570 67282 59600
rect 67398 59570 68066 59600
rect 68182 59570 68850 59600
rect 68966 59570 69634 59600
rect 69750 59570 70418 59600
rect 70534 59570 71202 59600
rect 71318 59570 71986 59600
rect 72102 59570 72770 59600
rect 72886 59570 73554 59600
rect 73670 59570 74338 59600
rect 74454 59570 75122 59600
rect 75238 59570 75906 59600
rect 76022 59570 76690 59600
rect 76806 59570 77474 59600
rect 77590 59570 78258 59600
rect 78374 59570 79042 59600
rect 79158 59570 79826 59600
rect 79942 59570 80610 59600
rect 80726 59570 81394 59600
rect 81510 59570 82178 59600
rect 82294 59570 82962 59600
rect 83078 59570 83746 59600
rect 83862 59570 84530 59600
rect 84646 59570 85314 59600
rect 85430 59570 86098 59600
rect 86214 59570 86882 59600
rect 86998 59570 87666 59600
rect 87782 59570 88450 59600
rect 88566 59570 89234 59600
rect 1470 430 89306 59570
rect 1470 400 3610 430
rect 3726 400 3778 430
rect 3894 400 3946 430
rect 4062 400 4114 430
rect 4230 400 4282 430
rect 4398 400 4450 430
rect 4566 400 4618 430
rect 4734 400 4786 430
rect 4902 400 4954 430
rect 5070 400 5122 430
rect 5238 400 5290 430
rect 5406 400 5458 430
rect 5574 400 5626 430
rect 5742 400 5794 430
rect 5910 400 5962 430
rect 6078 400 6130 430
rect 6246 400 6298 430
rect 6414 400 6466 430
rect 6582 400 6634 430
rect 6750 400 6802 430
rect 6918 400 6970 430
rect 7086 400 7138 430
rect 7254 400 7306 430
rect 7422 400 7474 430
rect 7590 400 7642 430
rect 7758 400 7810 430
rect 7926 400 7978 430
rect 8094 400 8146 430
rect 8262 400 8314 430
rect 8430 400 8482 430
rect 8598 400 8650 430
rect 8766 400 8818 430
rect 8934 400 8986 430
rect 9102 400 9154 430
rect 9270 400 9322 430
rect 9438 400 9490 430
rect 9606 400 9658 430
rect 9774 400 9826 430
rect 9942 400 9994 430
rect 10110 400 10162 430
rect 10278 400 10330 430
rect 10446 400 10498 430
rect 10614 400 10666 430
rect 10782 400 10834 430
rect 10950 400 11002 430
rect 11118 400 11170 430
rect 11286 400 11338 430
rect 11454 400 11506 430
rect 11622 400 11674 430
rect 11790 400 11842 430
rect 11958 400 12010 430
rect 12126 400 12178 430
rect 12294 400 12346 430
rect 12462 400 12514 430
rect 12630 400 12682 430
rect 12798 400 12850 430
rect 12966 400 13018 430
rect 13134 400 13186 430
rect 13302 400 13354 430
rect 13470 400 13522 430
rect 13638 400 13690 430
rect 13806 400 13858 430
rect 13974 400 14026 430
rect 14142 400 14194 430
rect 14310 400 14362 430
rect 14478 400 14530 430
rect 14646 400 14698 430
rect 14814 400 14866 430
rect 14982 400 15034 430
rect 15150 400 15202 430
rect 15318 400 15370 430
rect 15486 400 15538 430
rect 15654 400 15706 430
rect 15822 400 15874 430
rect 15990 400 16042 430
rect 16158 400 16210 430
rect 16326 400 16378 430
rect 16494 400 16546 430
rect 16662 400 16714 430
rect 16830 400 16882 430
rect 16998 400 17050 430
rect 17166 400 17218 430
rect 17334 400 17386 430
rect 17502 400 17554 430
rect 17670 400 17722 430
rect 17838 400 17890 430
rect 18006 400 18058 430
rect 18174 400 18226 430
rect 18342 400 18394 430
rect 18510 400 18562 430
rect 18678 400 18730 430
rect 18846 400 18898 430
rect 19014 400 19066 430
rect 19182 400 19234 430
rect 19350 400 19402 430
rect 19518 400 19570 430
rect 19686 400 19738 430
rect 19854 400 19906 430
rect 20022 400 20074 430
rect 20190 400 20242 430
rect 20358 400 20410 430
rect 20526 400 20578 430
rect 20694 400 20746 430
rect 20862 400 20914 430
rect 21030 400 21082 430
rect 21198 400 21250 430
rect 21366 400 21418 430
rect 21534 400 21586 430
rect 21702 400 21754 430
rect 21870 400 21922 430
rect 22038 400 22090 430
rect 22206 400 22258 430
rect 22374 400 22426 430
rect 22542 400 22594 430
rect 22710 400 22762 430
rect 22878 400 22930 430
rect 23046 400 23098 430
rect 23214 400 23266 430
rect 23382 400 23434 430
rect 23550 400 23602 430
rect 23718 400 23770 430
rect 23886 400 23938 430
rect 24054 400 24106 430
rect 24222 400 24274 430
rect 24390 400 24442 430
rect 24558 400 24610 430
rect 24726 400 24778 430
rect 24894 400 24946 430
rect 25062 400 25114 430
rect 25230 400 25282 430
rect 25398 400 25450 430
rect 25566 400 25618 430
rect 25734 400 25786 430
rect 25902 400 25954 430
rect 26070 400 26122 430
rect 26238 400 26290 430
rect 26406 400 26458 430
rect 26574 400 26626 430
rect 26742 400 26794 430
rect 26910 400 26962 430
rect 27078 400 27130 430
rect 27246 400 27298 430
rect 27414 400 27466 430
rect 27582 400 27634 430
rect 27750 400 27802 430
rect 27918 400 27970 430
rect 28086 400 28138 430
rect 28254 400 28306 430
rect 28422 400 28474 430
rect 28590 400 28642 430
rect 28758 400 28810 430
rect 28926 400 28978 430
rect 29094 400 29146 430
rect 29262 400 29314 430
rect 29430 400 29482 430
rect 29598 400 29650 430
rect 29766 400 29818 430
rect 29934 400 29986 430
rect 30102 400 30154 430
rect 30270 400 30322 430
rect 30438 400 30490 430
rect 30606 400 30658 430
rect 30774 400 30826 430
rect 30942 400 30994 430
rect 31110 400 31162 430
rect 31278 400 31330 430
rect 31446 400 31498 430
rect 31614 400 31666 430
rect 31782 400 31834 430
rect 31950 400 32002 430
rect 32118 400 32170 430
rect 32286 400 32338 430
rect 32454 400 32506 430
rect 32622 400 32674 430
rect 32790 400 32842 430
rect 32958 400 33010 430
rect 33126 400 33178 430
rect 33294 400 33346 430
rect 33462 400 33514 430
rect 33630 400 33682 430
rect 33798 400 33850 430
rect 33966 400 34018 430
rect 34134 400 34186 430
rect 34302 400 34354 430
rect 34470 400 34522 430
rect 34638 400 34690 430
rect 34806 400 34858 430
rect 34974 400 35026 430
rect 35142 400 35194 430
rect 35310 400 35362 430
rect 35478 400 35530 430
rect 35646 400 35698 430
rect 35814 400 35866 430
rect 35982 400 36034 430
rect 36150 400 36202 430
rect 36318 400 36370 430
rect 36486 400 36538 430
rect 36654 400 36706 430
rect 36822 400 36874 430
rect 36990 400 37042 430
rect 37158 400 37210 430
rect 37326 400 37378 430
rect 37494 400 37546 430
rect 37662 400 37714 430
rect 37830 400 37882 430
rect 37998 400 38050 430
rect 38166 400 38218 430
rect 38334 400 38386 430
rect 38502 400 38554 430
rect 38670 400 38722 430
rect 38838 400 38890 430
rect 39006 400 39058 430
rect 39174 400 39226 430
rect 39342 400 39394 430
rect 39510 400 39562 430
rect 39678 400 39730 430
rect 39846 400 39898 430
rect 40014 400 40066 430
rect 40182 400 40234 430
rect 40350 400 40402 430
rect 40518 400 40570 430
rect 40686 400 40738 430
rect 40854 400 40906 430
rect 41022 400 41074 430
rect 41190 400 41242 430
rect 41358 400 41410 430
rect 41526 400 41578 430
rect 41694 400 41746 430
rect 41862 400 41914 430
rect 42030 400 42082 430
rect 42198 400 42250 430
rect 42366 400 42418 430
rect 42534 400 42586 430
rect 42702 400 42754 430
rect 42870 400 42922 430
rect 43038 400 43090 430
rect 43206 400 43258 430
rect 43374 400 43426 430
rect 43542 400 43594 430
rect 43710 400 43762 430
rect 43878 400 43930 430
rect 44046 400 44098 430
rect 44214 400 44266 430
rect 44382 400 44434 430
rect 44550 400 44602 430
rect 44718 400 44770 430
rect 44886 400 44938 430
rect 45054 400 45106 430
rect 45222 400 45274 430
rect 45390 400 45442 430
rect 45558 400 45610 430
rect 45726 400 45778 430
rect 45894 400 45946 430
rect 46062 400 46114 430
rect 46230 400 46282 430
rect 46398 400 46450 430
rect 46566 400 46618 430
rect 46734 400 46786 430
rect 46902 400 46954 430
rect 47070 400 47122 430
rect 47238 400 47290 430
rect 47406 400 47458 430
rect 47574 400 47626 430
rect 47742 400 47794 430
rect 47910 400 47962 430
rect 48078 400 48130 430
rect 48246 400 48298 430
rect 48414 400 48466 430
rect 48582 400 48634 430
rect 48750 400 48802 430
rect 48918 400 48970 430
rect 49086 400 49138 430
rect 49254 400 49306 430
rect 49422 400 49474 430
rect 49590 400 49642 430
rect 49758 400 49810 430
rect 49926 400 49978 430
rect 50094 400 50146 430
rect 50262 400 50314 430
rect 50430 400 50482 430
rect 50598 400 50650 430
rect 50766 400 50818 430
rect 50934 400 50986 430
rect 51102 400 51154 430
rect 51270 400 51322 430
rect 51438 400 51490 430
rect 51606 400 51658 430
rect 51774 400 51826 430
rect 51942 400 51994 430
rect 52110 400 52162 430
rect 52278 400 52330 430
rect 52446 400 52498 430
rect 52614 400 52666 430
rect 52782 400 52834 430
rect 52950 400 53002 430
rect 53118 400 53170 430
rect 53286 400 53338 430
rect 53454 400 53506 430
rect 53622 400 53674 430
rect 53790 400 53842 430
rect 53958 400 54010 430
rect 54126 400 54178 430
rect 54294 400 54346 430
rect 54462 400 54514 430
rect 54630 400 54682 430
rect 54798 400 54850 430
rect 54966 400 55018 430
rect 55134 400 55186 430
rect 55302 400 55354 430
rect 55470 400 55522 430
rect 55638 400 55690 430
rect 55806 400 55858 430
rect 55974 400 56026 430
rect 56142 400 56194 430
rect 56310 400 56362 430
rect 56478 400 56530 430
rect 56646 400 56698 430
rect 56814 400 56866 430
rect 56982 400 57034 430
rect 57150 400 57202 430
rect 57318 400 57370 430
rect 57486 400 57538 430
rect 57654 400 57706 430
rect 57822 400 57874 430
rect 57990 400 58042 430
rect 58158 400 58210 430
rect 58326 400 58378 430
rect 58494 400 58546 430
rect 58662 400 58714 430
rect 58830 400 58882 430
rect 58998 400 59050 430
rect 59166 400 59218 430
rect 59334 400 59386 430
rect 59502 400 59554 430
rect 59670 400 59722 430
rect 59838 400 59890 430
rect 60006 400 60058 430
rect 60174 400 60226 430
rect 60342 400 60394 430
rect 60510 400 60562 430
rect 60678 400 60730 430
rect 60846 400 60898 430
rect 61014 400 61066 430
rect 61182 400 61234 430
rect 61350 400 61402 430
rect 61518 400 61570 430
rect 61686 400 61738 430
rect 61854 400 61906 430
rect 62022 400 62074 430
rect 62190 400 62242 430
rect 62358 400 62410 430
rect 62526 400 62578 430
rect 62694 400 62746 430
rect 62862 400 62914 430
rect 63030 400 63082 430
rect 63198 400 63250 430
rect 63366 400 63418 430
rect 63534 400 63586 430
rect 63702 400 63754 430
rect 63870 400 63922 430
rect 64038 400 64090 430
rect 64206 400 64258 430
rect 64374 400 64426 430
rect 64542 400 64594 430
rect 64710 400 64762 430
rect 64878 400 64930 430
rect 65046 400 65098 430
rect 65214 400 65266 430
rect 65382 400 65434 430
rect 65550 400 65602 430
rect 65718 400 65770 430
rect 65886 400 65938 430
rect 66054 400 66106 430
rect 66222 400 66274 430
rect 66390 400 66442 430
rect 66558 400 66610 430
rect 66726 400 66778 430
rect 66894 400 66946 430
rect 67062 400 67114 430
rect 67230 400 67282 430
rect 67398 400 67450 430
rect 67566 400 67618 430
rect 67734 400 67786 430
rect 67902 400 67954 430
rect 68070 400 68122 430
rect 68238 400 68290 430
rect 68406 400 68458 430
rect 68574 400 68626 430
rect 68742 400 68794 430
rect 68910 400 68962 430
rect 69078 400 69130 430
rect 69246 400 69298 430
rect 69414 400 69466 430
rect 69582 400 69634 430
rect 69750 400 69802 430
rect 69918 400 69970 430
rect 70086 400 70138 430
rect 70254 400 70306 430
rect 70422 400 70474 430
rect 70590 400 70642 430
rect 70758 400 70810 430
rect 70926 400 70978 430
rect 71094 400 71146 430
rect 71262 400 71314 430
rect 71430 400 71482 430
rect 71598 400 71650 430
rect 71766 400 71818 430
rect 71934 400 71986 430
rect 72102 400 72154 430
rect 72270 400 72322 430
rect 72438 400 72490 430
rect 72606 400 72658 430
rect 72774 400 72826 430
rect 72942 400 72994 430
rect 73110 400 73162 430
rect 73278 400 73330 430
rect 73446 400 73498 430
rect 73614 400 73666 430
rect 73782 400 73834 430
rect 73950 400 74002 430
rect 74118 400 74170 430
rect 74286 400 74338 430
rect 74454 400 74506 430
rect 74622 400 74674 430
rect 74790 400 74842 430
rect 74958 400 75010 430
rect 75126 400 75178 430
rect 75294 400 75346 430
rect 75462 400 75514 430
rect 75630 400 75682 430
rect 75798 400 75850 430
rect 75966 400 76018 430
rect 76134 400 76186 430
rect 76302 400 76354 430
rect 76470 400 76522 430
rect 76638 400 76690 430
rect 76806 400 76858 430
rect 76974 400 77026 430
rect 77142 400 77194 430
rect 77310 400 77362 430
rect 77478 400 77530 430
rect 77646 400 77698 430
rect 77814 400 77866 430
rect 77982 400 78034 430
rect 78150 400 78202 430
rect 78318 400 78370 430
rect 78486 400 78538 430
rect 78654 400 78706 430
rect 78822 400 78874 430
rect 78990 400 79042 430
rect 79158 400 79210 430
rect 79326 400 79378 430
rect 79494 400 79546 430
rect 79662 400 79714 430
rect 79830 400 79882 430
rect 79998 400 80050 430
rect 80166 400 80218 430
rect 80334 400 80386 430
rect 80502 400 80554 430
rect 80670 400 80722 430
rect 80838 400 80890 430
rect 81006 400 81058 430
rect 81174 400 81226 430
rect 81342 400 81394 430
rect 81510 400 81562 430
rect 81678 400 81730 430
rect 81846 400 81898 430
rect 82014 400 82066 430
rect 82182 400 82234 430
rect 82350 400 82402 430
rect 82518 400 82570 430
rect 82686 400 82738 430
rect 82854 400 82906 430
rect 83022 400 83074 430
rect 83190 400 83242 430
rect 83358 400 83410 430
rect 83526 400 83578 430
rect 83694 400 83746 430
rect 83862 400 83914 430
rect 84030 400 84082 430
rect 84198 400 84250 430
rect 84366 400 84418 430
rect 84534 400 84586 430
rect 84702 400 84754 430
rect 84870 400 84922 430
rect 85038 400 85090 430
rect 85206 400 85258 430
rect 85374 400 85426 430
rect 85542 400 85594 430
rect 85710 400 85762 430
rect 85878 400 85930 430
rect 86046 400 86098 430
rect 86214 400 86266 430
rect 86382 400 89306 430
<< obsm3 >>
rect 1465 406 89311 58786
<< metal4 >>
rect 2224 1538 2384 58438
rect 9904 1538 10064 58438
rect 17584 1538 17744 58438
rect 25264 1538 25424 58438
rect 32944 1538 33104 58438
rect 40624 1538 40784 58438
rect 48304 1538 48464 58438
rect 55984 1538 56144 58438
rect 63664 1538 63824 58438
rect 71344 1538 71504 58438
rect 79024 1538 79184 58438
rect 86704 1538 86864 58438
<< obsm4 >>
rect 8526 1508 9874 58119
rect 10094 1508 17554 58119
rect 17774 1508 25234 58119
rect 25454 1508 32914 58119
rect 33134 1508 40594 58119
rect 40814 1508 48274 58119
rect 48494 1508 49378 58119
rect 8526 625 49378 1508
<< labels >>
rlabel metal2 s 672 59600 728 60000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 24192 59600 24248 60000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 26544 59600 26600 60000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 28896 59600 28952 60000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 31248 59600 31304 60000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 33600 59600 33656 60000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 35952 59600 36008 60000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 38304 59600 38360 60000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 40656 59600 40712 60000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 43008 59600 43064 60000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 45360 59600 45416 60000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3024 59600 3080 60000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 47712 59600 47768 60000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 50064 59600 50120 60000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 52416 59600 52472 60000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 54768 59600 54824 60000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 57120 59600 57176 60000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 59472 59600 59528 60000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 61824 59600 61880 60000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 64176 59600 64232 60000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 66528 59600 66584 60000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 68880 59600 68936 60000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 5376 59600 5432 60000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 71232 59600 71288 60000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 73584 59600 73640 60000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 75936 59600 75992 60000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 78288 59600 78344 60000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 80640 59600 80696 60000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 82992 59600 83048 60000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 85344 59600 85400 60000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 87696 59600 87752 60000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 7728 59600 7784 60000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 10080 59600 10136 60000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 12432 59600 12488 60000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 14784 59600 14840 60000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 17136 59600 17192 60000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 19488 59600 19544 60000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 21840 59600 21896 60000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1456 59600 1512 60000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 24976 59600 25032 60000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 27328 59600 27384 60000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 29680 59600 29736 60000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 32032 59600 32088 60000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 34384 59600 34440 60000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 36736 59600 36792 60000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 39088 59600 39144 60000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 41440 59600 41496 60000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 43792 59600 43848 60000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 46144 59600 46200 60000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 3808 59600 3864 60000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 48496 59600 48552 60000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 50848 59600 50904 60000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 53200 59600 53256 60000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 55552 59600 55608 60000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 57904 59600 57960 60000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 60256 59600 60312 60000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 62608 59600 62664 60000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 64960 59600 65016 60000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 67312 59600 67368 60000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 69664 59600 69720 60000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 6160 59600 6216 60000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 72016 59600 72072 60000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 74368 59600 74424 60000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 76720 59600 76776 60000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 79072 59600 79128 60000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 81424 59600 81480 60000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 83776 59600 83832 60000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 86128 59600 86184 60000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 88480 59600 88536 60000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 8512 59600 8568 60000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 10864 59600 10920 60000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 13216 59600 13272 60000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 15568 59600 15624 60000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 17920 59600 17976 60000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 20272 59600 20328 60000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 22624 59600 22680 60000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2240 59600 2296 60000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 25760 59600 25816 60000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 28112 59600 28168 60000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 30464 59600 30520 60000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 32816 59600 32872 60000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 35168 59600 35224 60000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 37520 59600 37576 60000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 39872 59600 39928 60000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 42224 59600 42280 60000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 44576 59600 44632 60000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 46928 59600 46984 60000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 4592 59600 4648 60000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 49280 59600 49336 60000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 51632 59600 51688 60000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 53984 59600 54040 60000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 56336 59600 56392 60000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 58688 59600 58744 60000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 61040 59600 61096 60000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 63392 59600 63448 60000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 65744 59600 65800 60000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 68096 59600 68152 60000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 70448 59600 70504 60000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 6944 59600 7000 60000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 72800 59600 72856 60000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 75152 59600 75208 60000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 77504 59600 77560 60000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 79856 59600 79912 60000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 82208 59600 82264 60000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 84560 59600 84616 60000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 86912 59600 86968 60000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 89264 59600 89320 60000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 9296 59600 9352 60000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 11648 59600 11704 60000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 14000 59600 14056 60000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 16352 59600 16408 60000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 18704 59600 18760 60000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 21056 59600 21112 60000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 23408 59600 23464 60000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 85960 0 86016 400 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 86128 0 86184 400 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 86296 0 86352 400 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 21448 0 21504 400 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 71848 0 71904 400 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 72856 0 72912 400 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 73360 0 73416 400 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 73864 0 73920 400 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 74368 0 74424 400 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 74872 0 74928 400 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 75376 0 75432 400 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 75880 0 75936 400 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 26488 0 26544 400 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 76888 0 76944 400 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 77392 0 77448 400 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 77896 0 77952 400 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 78400 0 78456 400 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 78904 0 78960 400 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 79912 0 79968 400 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 80920 0 80976 400 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 81424 0 81480 400 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 81928 0 81984 400 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 82432 0 82488 400 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 82936 0 82992 400 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 83944 0 84000 400 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 84952 0 85008 400 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 85456 0 85512 400 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 27496 0 27552 400 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 28504 0 28560 400 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 29008 0 29064 400 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 29512 0 29568 400 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 30520 0 30576 400 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 21952 0 22008 400 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 31528 0 31584 400 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 32536 0 32592 400 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 33040 0 33096 400 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 33544 0 33600 400 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 34552 0 34608 400 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 35056 0 35112 400 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 35560 0 35616 400 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 36064 0 36120 400 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 22456 0 22512 400 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 36568 0 36624 400 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 37072 0 37128 400 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 37576 0 37632 400 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 38080 0 38136 400 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 38584 0 38640 400 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 39592 0 39648 400 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 40600 0 40656 400 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 22960 0 23016 400 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 41608 0 41664 400 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 42616 0 42672 400 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 43120 0 43176 400 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 43624 0 43680 400 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 44632 0 44688 400 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 45136 0 45192 400 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 45640 0 45696 400 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 46144 0 46200 400 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 23464 0 23520 400 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 46648 0 46704 400 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 47656 0 47712 400 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 48664 0 48720 400 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 49168 0 49224 400 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 49672 0 49728 400 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 50176 0 50232 400 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 50680 0 50736 400 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 51184 0 51240 400 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 51688 0 51744 400 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 52192 0 52248 400 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 52696 0 52752 400 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 53200 0 53256 400 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 53704 0 53760 400 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 54208 0 54264 400 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 54712 0 54768 400 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 55720 0 55776 400 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 24472 0 24528 400 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 56728 0 56784 400 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 57232 0 57288 400 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 57736 0 57792 400 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 58240 0 58296 400 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 58744 0 58800 400 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 59248 0 59304 400 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 59752 0 59808 400 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 60256 0 60312 400 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 60760 0 60816 400 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 61264 0 61320 400 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 24976 0 25032 400 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 61768 0 61824 400 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 62272 0 62328 400 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 62776 0 62832 400 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 63784 0 63840 400 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 64792 0 64848 400 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 65296 0 65352 400 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 65800 0 65856 400 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 66304 0 66360 400 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 25480 0 25536 400 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 66808 0 66864 400 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 67312 0 67368 400 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 67816 0 67872 400 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 68824 0 68880 400 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 69832 0 69888 400 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 70840 0 70896 400 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 72016 0 72072 400 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 72520 0 72576 400 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 73024 0 73080 400 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 73528 0 73584 400 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 74032 0 74088 400 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 74536 0 74592 400 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 75040 0 75096 400 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 75544 0 75600 400 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 76048 0 76104 400 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 76552 0 76608 400 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 26656 0 26712 400 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 77056 0 77112 400 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 77560 0 77616 400 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 78064 0 78120 400 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 78568 0 78624 400 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 79072 0 79128 400 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 79576 0 79632 400 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 80080 0 80136 400 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 80584 0 80640 400 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 81088 0 81144 400 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 81592 0 81648 400 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 27160 0 27216 400 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 82096 0 82152 400 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 82600 0 82656 400 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 83104 0 83160 400 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 83608 0 83664 400 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 84112 0 84168 400 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 84616 0 84672 400 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 85120 0 85176 400 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 85624 0 85680 400 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 27664 0 27720 400 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 28168 0 28224 400 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 29176 0 29232 400 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 30184 0 30240 400 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 31192 0 31248 400 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 22120 0 22176 400 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 31696 0 31752 400 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 32200 0 32256 400 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 32704 0 32760 400 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 33208 0 33264 400 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 33712 0 33768 400 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 34216 0 34272 400 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 34720 0 34776 400 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 35224 0 35280 400 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 35728 0 35784 400 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 36232 0 36288 400 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 22624 0 22680 400 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 36736 0 36792 400 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 37240 0 37296 400 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 37744 0 37800 400 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 38248 0 38304 400 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 38752 0 38808 400 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 39256 0 39312 400 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 39760 0 39816 400 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 40264 0 40320 400 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 40768 0 40824 400 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 41272 0 41328 400 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 23128 0 23184 400 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 41776 0 41832 400 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 42280 0 42336 400 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 42784 0 42840 400 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 43288 0 43344 400 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 43792 0 43848 400 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 44296 0 44352 400 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 44800 0 44856 400 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 45304 0 45360 400 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 45808 0 45864 400 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 46312 0 46368 400 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 23632 0 23688 400 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 46816 0 46872 400 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 47320 0 47376 400 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 47824 0 47880 400 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 48328 0 48384 400 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 48832 0 48888 400 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 49336 0 49392 400 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 49840 0 49896 400 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 50344 0 50400 400 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 50848 0 50904 400 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 51352 0 51408 400 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 24136 0 24192 400 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 51856 0 51912 400 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 52360 0 52416 400 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 52864 0 52920 400 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 53368 0 53424 400 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 53872 0 53928 400 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 54376 0 54432 400 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 54880 0 54936 400 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 55384 0 55440 400 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 55888 0 55944 400 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 56392 0 56448 400 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 24640 0 24696 400 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 56896 0 56952 400 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 57400 0 57456 400 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 57904 0 57960 400 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 58408 0 58464 400 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 58912 0 58968 400 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 59416 0 59472 400 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 59920 0 59976 400 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 60424 0 60480 400 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 60928 0 60984 400 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 61432 0 61488 400 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 25144 0 25200 400 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 62440 0 62496 400 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 62944 0 63000 400 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 63448 0 63504 400 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 63952 0 64008 400 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 64456 0 64512 400 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 64960 0 65016 400 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 65464 0 65520 400 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 65968 0 66024 400 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 66472 0 66528 400 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 25648 0 25704 400 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 66976 0 67032 400 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 67480 0 67536 400 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 67984 0 68040 400 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 68488 0 68544 400 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 68992 0 69048 400 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 69496 0 69552 400 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 70000 0 70056 400 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 70504 0 70560 400 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 71008 0 71064 400 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 71512 0 71568 400 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 26152 0 26208 400 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 21784 0 21840 400 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 72184 0 72240 400 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 72688 0 72744 400 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 73192 0 73248 400 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 73696 0 73752 400 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 74200 0 74256 400 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 74704 0 74760 400 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 75208 0 75264 400 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 75712 0 75768 400 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 76216 0 76272 400 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 26824 0 26880 400 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 77224 0 77280 400 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 78232 0 78288 400 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 78736 0 78792 400 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 79240 0 79296 400 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 79744 0 79800 400 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 80248 0 80304 400 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 80752 0 80808 400 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 81256 0 81312 400 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 81760 0 81816 400 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 82264 0 82320 400 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 82768 0 82824 400 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 83272 0 83328 400 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 83776 0 83832 400 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 84280 0 84336 400 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 85288 0 85344 400 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 85792 0 85848 400 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 27832 0 27888 400 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 28840 0 28896 400 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 29848 0 29904 400 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 30352 0 30408 400 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 30856 0 30912 400 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 31864 0 31920 400 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 32368 0 32424 400 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 32872 0 32928 400 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 33880 0 33936 400 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 34384 0 34440 400 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 34888 0 34944 400 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 35896 0 35952 400 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 22792 0 22848 400 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 36904 0 36960 400 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 37912 0 37968 400 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 38416 0 38472 400 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 38920 0 38976 400 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 39928 0 39984 400 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 40432 0 40488 400 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 40936 0 40992 400 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 41440 0 41496 400 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 41944 0 42000 400 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 42448 0 42504 400 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 42952 0 43008 400 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 43456 0 43512 400 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 43960 0 44016 400 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 44968 0 45024 400 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 45976 0 46032 400 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 46480 0 46536 400 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 23800 0 23856 400 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 46984 0 47040 400 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 47488 0 47544 400 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 47992 0 48048 400 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 48496 0 48552 400 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 49000 0 49056 400 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 50008 0 50064 400 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 51016 0 51072 400 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 52024 0 52080 400 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 53032 0 53088 400 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 54040 0 54096 400 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 54544 0 54600 400 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 55048 0 55104 400 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 55552 0 55608 400 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 56056 0 56112 400 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 56560 0 56616 400 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 24808 0 24864 400 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 57064 0 57120 400 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 57568 0 57624 400 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 58072 0 58128 400 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 58576 0 58632 400 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 59080 0 59136 400 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 59584 0 59640 400 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 60088 0 60144 400 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 60592 0 60648 400 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 61096 0 61152 400 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 62104 0 62160 400 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 62608 0 62664 400 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 63112 0 63168 400 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 63616 0 63672 400 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 64120 0 64176 400 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 65128 0 65184 400 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 65632 0 65688 400 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 66136 0 66192 400 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 66640 0 66696 400 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 25816 0 25872 400 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 67144 0 67200 400 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 68152 0 68208 400 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 69160 0 69216 400 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 70168 0 70224 400 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 70672 0 70728 400 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 71176 0 71232 400 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 71680 0 71736 400 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 26320 0 26376 400 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 2224 1538 2384 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 58438 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 58438 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 3640 0 3696 400 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 3808 0 3864 400 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 3976 0 4032 400 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 4648 0 4704 400 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 10360 0 10416 400 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 11368 0 11424 400 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 12376 0 12432 400 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 13384 0 13440 400 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 14392 0 14448 400 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 5320 0 5376 400 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 15400 0 15456 400 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 16408 0 16464 400 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 16912 0 16968 400 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 17416 0 17472 400 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 18424 0 18480 400 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 19432 0 19488 400 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 19936 0 19992 400 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 5992 0 6048 400 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 20440 0 20496 400 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 20944 0 21000 400 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 6664 0 6720 400 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 7336 0 7392 400 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 7840 0 7896 400 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 8344 0 8400 400 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 8848 0 8904 400 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 9352 0 9408 400 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 9856 0 9912 400 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 4144 0 4200 400 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 4816 0 4872 400 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 11032 0 11088 400 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 11536 0 11592 400 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 12040 0 12096 400 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 12544 0 12600 400 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 13048 0 13104 400 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 13552 0 13608 400 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 14056 0 14112 400 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 15064 0 15120 400 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 5488 0 5544 400 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 15568 0 15624 400 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 16072 0 16128 400 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 17080 0 17136 400 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 18088 0 18144 400 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 19096 0 19152 400 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 19600 0 19656 400 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 20104 0 20160 400 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 6160 0 6216 400 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 20608 0 20664 400 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 21112 0 21168 400 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 6832 0 6888 400 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 7504 0 7560 400 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 8008 0 8064 400 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 8512 0 8568 400 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 9016 0 9072 400 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 10024 0 10080 400 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 4984 0 5040 400 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 10696 0 10752 400 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 11200 0 11256 400 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 11704 0 11760 400 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 12208 0 12264 400 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 12712 0 12768 400 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 13216 0 13272 400 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 13720 0 13776 400 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 14224 0 14280 400 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 14728 0 14784 400 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 5656 0 5712 400 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 15736 0 15792 400 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 16744 0 16800 400 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 17752 0 17808 400 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 18256 0 18312 400 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 18760 0 18816 400 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 19264 0 19320 400 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 19768 0 19824 400 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 20272 0 20328 400 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 6328 0 6384 400 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 20776 0 20832 400 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 21280 0 21336 400 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 7000 0 7056 400 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 7672 0 7728 400 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 8176 0 8232 400 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 8680 0 8736 400 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 9184 0 9240 400 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 9688 0 9744 400 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 10192 0 10248 400 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 5152 0 5208 400 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 5824 0 5880 400 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 6496 0 6552 400 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 7168 0 7224 400 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 4312 0 4368 400 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 4480 0 4536 400 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 90000 60000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3593948
string GDS_FILE /Volumes/Efabless/ParaRAM/openlane/user_proj_example/runs/22_11_05_15_51/results/signoff/user_proj_example.magic.gds
string GDS_START 205212
<< end >>

