magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -81 602 81 608
rect -81 576 -75 602
rect -49 576 -13 602
rect 13 576 49 602
rect 75 576 81 602
rect -81 540 81 576
rect -81 514 -75 540
rect -49 514 -13 540
rect 13 514 49 540
rect 75 514 81 540
rect -81 478 81 514
rect -81 452 -75 478
rect -49 452 -13 478
rect 13 452 49 478
rect 75 452 81 478
rect -81 416 81 452
rect -81 390 -75 416
rect -49 390 -13 416
rect 13 390 49 416
rect 75 390 81 416
rect -81 354 81 390
rect -81 328 -75 354
rect -49 328 -13 354
rect 13 328 49 354
rect 75 328 81 354
rect -81 292 81 328
rect -81 266 -75 292
rect -49 266 -13 292
rect 13 266 49 292
rect 75 266 81 292
rect -81 230 81 266
rect -81 204 -75 230
rect -49 204 -13 230
rect 13 204 49 230
rect 75 204 81 230
rect -81 168 81 204
rect -81 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 81 168
rect -81 106 81 142
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -142 81 -106
rect -81 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 81 -142
rect -81 -204 81 -168
rect -81 -230 -75 -204
rect -49 -230 -13 -204
rect 13 -230 49 -204
rect 75 -230 81 -204
rect -81 -266 81 -230
rect -81 -292 -75 -266
rect -49 -292 -13 -266
rect 13 -292 49 -266
rect 75 -292 81 -266
rect -81 -328 81 -292
rect -81 -354 -75 -328
rect -49 -354 -13 -328
rect 13 -354 49 -328
rect 75 -354 81 -328
rect -81 -390 81 -354
rect -81 -416 -75 -390
rect -49 -416 -13 -390
rect 13 -416 49 -390
rect 75 -416 81 -390
rect -81 -452 81 -416
rect -81 -478 -75 -452
rect -49 -478 -13 -452
rect 13 -478 49 -452
rect 75 -478 81 -452
rect -81 -514 81 -478
rect -81 -540 -75 -514
rect -49 -540 -13 -514
rect 13 -540 49 -514
rect 75 -540 81 -514
rect -81 -576 81 -540
rect -81 -602 -75 -576
rect -49 -602 -13 -576
rect 13 -602 49 -576
rect 75 -602 81 -576
rect -81 -608 81 -602
<< via1 >>
rect -75 576 -49 602
rect -13 576 13 602
rect 49 576 75 602
rect -75 514 -49 540
rect -13 514 13 540
rect 49 514 75 540
rect -75 452 -49 478
rect -13 452 13 478
rect 49 452 75 478
rect -75 390 -49 416
rect -13 390 13 416
rect 49 390 75 416
rect -75 328 -49 354
rect -13 328 13 354
rect 49 328 75 354
rect -75 266 -49 292
rect -13 266 13 292
rect 49 266 75 292
rect -75 204 -49 230
rect -13 204 13 230
rect 49 204 75 230
rect -75 142 -49 168
rect -13 142 13 168
rect 49 142 75 168
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
rect -75 -168 -49 -142
rect -13 -168 13 -142
rect 49 -168 75 -142
rect -75 -230 -49 -204
rect -13 -230 13 -204
rect 49 -230 75 -204
rect -75 -292 -49 -266
rect -13 -292 13 -266
rect 49 -292 75 -266
rect -75 -354 -49 -328
rect -13 -354 13 -328
rect 49 -354 75 -328
rect -75 -416 -49 -390
rect -13 -416 13 -390
rect 49 -416 75 -390
rect -75 -478 -49 -452
rect -13 -478 13 -452
rect 49 -478 75 -452
rect -75 -540 -49 -514
rect -13 -540 13 -514
rect 49 -540 75 -514
rect -75 -602 -49 -576
rect -13 -602 13 -576
rect 49 -602 75 -576
<< metal2 >>
rect -81 602 81 608
rect -81 576 -75 602
rect -49 576 -13 602
rect 13 576 49 602
rect 75 576 81 602
rect -81 540 81 576
rect -81 514 -75 540
rect -49 514 -13 540
rect 13 514 49 540
rect 75 514 81 540
rect -81 478 81 514
rect -81 452 -75 478
rect -49 452 -13 478
rect 13 452 49 478
rect 75 452 81 478
rect -81 416 81 452
rect -81 390 -75 416
rect -49 390 -13 416
rect 13 390 49 416
rect 75 390 81 416
rect -81 354 81 390
rect -81 328 -75 354
rect -49 328 -13 354
rect 13 328 49 354
rect 75 328 81 354
rect -81 292 81 328
rect -81 266 -75 292
rect -49 266 -13 292
rect 13 266 49 292
rect 75 266 81 292
rect -81 230 81 266
rect -81 204 -75 230
rect -49 204 -13 230
rect 13 204 49 230
rect 75 204 81 230
rect -81 168 81 204
rect -81 142 -75 168
rect -49 142 -13 168
rect 13 142 49 168
rect 75 142 81 168
rect -81 106 81 142
rect -81 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 81 106
rect -81 44 81 80
rect -81 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 81 44
rect -81 -18 81 18
rect -81 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 81 -18
rect -81 -80 81 -44
rect -81 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 81 -80
rect -81 -142 81 -106
rect -81 -168 -75 -142
rect -49 -168 -13 -142
rect 13 -168 49 -142
rect 75 -168 81 -142
rect -81 -204 81 -168
rect -81 -230 -75 -204
rect -49 -230 -13 -204
rect 13 -230 49 -204
rect 75 -230 81 -204
rect -81 -266 81 -230
rect -81 -292 -75 -266
rect -49 -292 -13 -266
rect 13 -292 49 -266
rect 75 -292 81 -266
rect -81 -328 81 -292
rect -81 -354 -75 -328
rect -49 -354 -13 -328
rect 13 -354 49 -328
rect 75 -354 81 -328
rect -81 -390 81 -354
rect -81 -416 -75 -390
rect -49 -416 -13 -390
rect 13 -416 49 -390
rect 75 -416 81 -390
rect -81 -452 81 -416
rect -81 -478 -75 -452
rect -49 -478 -13 -452
rect 13 -478 49 -452
rect 75 -478 81 -452
rect -81 -514 81 -478
rect -81 -540 -75 -514
rect -49 -540 -13 -514
rect 13 -540 49 -514
rect 75 -540 81 -514
rect -81 -576 81 -540
rect -81 -602 -75 -576
rect -49 -602 -13 -576
rect 13 -602 49 -576
rect 75 -602 81 -576
rect -81 -608 81 -602
<< properties >>
string GDS_END 1481186
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1477214
<< end >>
