magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -19 355 19 360
rect -19 327 -14 355
rect 14 327 19 355
rect -19 293 19 327
rect -19 265 -14 293
rect 14 265 19 293
rect -19 231 19 265
rect -19 203 -14 231
rect 14 203 19 231
rect -19 169 19 203
rect -19 141 -14 169
rect 14 141 19 169
rect -19 107 19 141
rect -19 79 -14 107
rect 14 79 19 107
rect -19 45 19 79
rect -19 17 -14 45
rect 14 17 19 45
rect -19 -17 19 17
rect -19 -45 -14 -17
rect 14 -45 19 -17
rect -19 -79 19 -45
rect -19 -107 -14 -79
rect 14 -107 19 -79
rect -19 -141 19 -107
rect -19 -169 -14 -141
rect 14 -169 19 -141
rect -19 -203 19 -169
rect -19 -231 -14 -203
rect 14 -231 19 -203
rect -19 -265 19 -231
rect -19 -293 -14 -265
rect 14 -293 19 -265
rect -19 -327 19 -293
rect -19 -355 -14 -327
rect 14 -355 19 -327
rect -19 -360 19 -355
<< via2 >>
rect -14 327 14 355
rect -14 265 14 293
rect -14 203 14 231
rect -14 141 14 169
rect -14 79 14 107
rect -14 17 14 45
rect -14 -45 14 -17
rect -14 -107 14 -79
rect -14 -169 14 -141
rect -14 -231 14 -203
rect -14 -293 14 -265
rect -14 -355 14 -327
<< metal3 >>
rect -19 355 19 360
rect -19 327 -14 355
rect 14 327 19 355
rect -19 293 19 327
rect -19 265 -14 293
rect 14 265 19 293
rect -19 231 19 265
rect -19 203 -14 231
rect 14 203 19 231
rect -19 169 19 203
rect -19 141 -14 169
rect 14 141 19 169
rect -19 107 19 141
rect -19 79 -14 107
rect 14 79 19 107
rect -19 45 19 79
rect -19 17 -14 45
rect 14 17 19 45
rect -19 -17 19 17
rect -19 -45 -14 -17
rect 14 -45 19 -17
rect -19 -79 19 -45
rect -19 -107 -14 -79
rect 14 -107 19 -79
rect -19 -141 19 -107
rect -19 -169 -14 -141
rect 14 -169 19 -141
rect -19 -203 19 -169
rect -19 -231 -14 -203
rect 14 -231 19 -203
rect -19 -265 19 -231
rect -19 -293 -14 -265
rect 14 -293 19 -265
rect -19 -327 19 -293
rect -19 -355 -14 -327
rect 14 -355 19 -327
rect -19 -360 19 -355
<< properties >>
string GDS_END 617514
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 616614
<< end >>
