magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 4006 1094
<< pwell >>
rect -86 -86 4006 453
<< mvnmos >>
rect 124 69 244 333
rect 348 69 468 333
rect 572 69 692 333
rect 796 69 916 333
rect 1020 69 1140 333
rect 1244 69 1364 333
rect 1468 69 1588 333
rect 1692 69 1812 333
rect 1916 69 2036 333
rect 2140 69 2260 333
rect 2364 69 2484 333
rect 2588 69 2708 333
rect 2916 69 3036 333
rect 3140 69 3260 333
rect 3364 69 3484 333
rect 3588 69 3708 333
<< mvpmos >>
rect 144 573 244 939
rect 368 573 468 939
rect 582 573 682 939
rect 806 573 906 939
rect 1030 573 1130 939
rect 1254 573 1354 939
rect 1478 573 1578 939
rect 1712 573 1812 939
rect 1926 573 2026 939
rect 2150 573 2250 939
rect 2374 573 2474 939
rect 2588 573 2688 939
rect 2936 610 3036 939
rect 3170 610 3270 939
rect 3374 610 3474 939
rect 3598 610 3698 939
<< mvndiff >>
rect 36 312 124 333
rect 36 172 49 312
rect 95 172 124 312
rect 36 69 124 172
rect 244 285 348 333
rect 244 239 273 285
rect 319 239 348 285
rect 244 69 348 239
rect 468 218 572 333
rect 468 172 497 218
rect 543 172 572 218
rect 468 69 572 172
rect 692 274 796 333
rect 692 228 721 274
rect 767 228 796 274
rect 692 69 796 228
rect 916 218 1020 333
rect 916 172 945 218
rect 991 172 1020 218
rect 916 69 1020 172
rect 1140 274 1244 333
rect 1140 228 1169 274
rect 1215 228 1244 274
rect 1140 69 1244 228
rect 1364 218 1468 333
rect 1364 172 1393 218
rect 1439 172 1468 218
rect 1364 69 1468 172
rect 1588 274 1692 333
rect 1588 228 1617 274
rect 1663 228 1692 274
rect 1588 69 1692 228
rect 1812 216 1916 333
rect 1812 170 1841 216
rect 1887 170 1916 216
rect 1812 69 1916 170
rect 2036 274 2140 333
rect 2036 228 2065 274
rect 2111 228 2140 274
rect 2036 69 2140 228
rect 2260 294 2364 333
rect 2260 154 2289 294
rect 2335 154 2364 294
rect 2260 69 2364 154
rect 2484 285 2588 333
rect 2484 239 2513 285
rect 2559 239 2588 285
rect 2484 69 2588 239
rect 2708 312 2916 333
rect 2708 172 2785 312
rect 2831 172 2916 312
rect 2708 69 2916 172
rect 3036 305 3140 333
rect 3036 165 3065 305
rect 3111 165 3140 305
rect 3036 69 3140 165
rect 3260 312 3364 333
rect 3260 172 3289 312
rect 3335 172 3364 312
rect 3260 69 3364 172
rect 3484 305 3588 333
rect 3484 165 3513 305
rect 3559 165 3588 305
rect 3484 69 3588 165
rect 3708 312 3796 333
rect 3708 172 3737 312
rect 3783 172 3796 312
rect 3708 69 3796 172
<< mvpdiff >>
rect 56 861 144 939
rect 56 721 69 861
rect 115 721 144 861
rect 56 573 144 721
rect 244 861 368 939
rect 244 721 273 861
rect 319 721 368 861
rect 244 573 368 721
rect 468 861 582 939
rect 468 721 497 861
rect 543 721 582 861
rect 468 573 582 721
rect 682 861 806 939
rect 682 721 711 861
rect 757 721 806 861
rect 682 573 806 721
rect 906 573 1030 939
rect 1130 573 1254 939
rect 1354 767 1478 939
rect 1354 721 1403 767
rect 1449 721 1478 767
rect 1354 573 1478 721
rect 1578 573 1712 939
rect 1812 870 1926 939
rect 1812 824 1841 870
rect 1887 824 1926 870
rect 1812 573 1926 824
rect 2026 573 2150 939
rect 2250 767 2374 939
rect 2250 721 2279 767
rect 2325 721 2374 767
rect 2250 573 2374 721
rect 2474 573 2588 939
rect 2688 870 2776 939
rect 2688 824 2717 870
rect 2763 824 2776 870
rect 2688 573 2776 824
rect 2848 926 2936 939
rect 2848 786 2861 926
rect 2907 786 2936 926
rect 2848 610 2936 786
rect 3036 861 3170 939
rect 3036 721 3065 861
rect 3111 721 3170 861
rect 3036 610 3170 721
rect 3270 861 3374 939
rect 3270 721 3299 861
rect 3345 721 3374 861
rect 3270 610 3374 721
rect 3474 861 3598 939
rect 3474 721 3503 861
rect 3549 721 3598 861
rect 3474 610 3598 721
rect 3698 861 3786 939
rect 3698 721 3727 861
rect 3773 721 3786 861
rect 3698 610 3786 721
<< mvndiffc >>
rect 49 172 95 312
rect 273 239 319 285
rect 497 172 543 218
rect 721 228 767 274
rect 945 172 991 218
rect 1169 228 1215 274
rect 1393 172 1439 218
rect 1617 228 1663 274
rect 1841 170 1887 216
rect 2065 228 2111 274
rect 2289 154 2335 294
rect 2513 239 2559 285
rect 2785 172 2831 312
rect 3065 165 3111 305
rect 3289 172 3335 312
rect 3513 165 3559 305
rect 3737 172 3783 312
<< mvpdiffc >>
rect 69 721 115 861
rect 273 721 319 861
rect 497 721 543 861
rect 711 721 757 861
rect 1403 721 1449 767
rect 1841 824 1887 870
rect 2279 721 2325 767
rect 2717 824 2763 870
rect 2861 786 2907 926
rect 3065 721 3111 861
rect 3299 721 3345 861
rect 3503 721 3549 861
rect 3727 721 3773 861
<< polysilicon >>
rect 144 939 244 983
rect 368 939 468 983
rect 582 939 682 983
rect 806 939 906 983
rect 1030 939 1130 983
rect 1254 939 1354 983
rect 1478 939 1578 983
rect 1712 939 1812 983
rect 1926 939 2026 983
rect 2150 939 2250 983
rect 2374 939 2474 983
rect 2588 939 2688 983
rect 2936 939 3036 983
rect 3170 939 3270 983
rect 3374 939 3474 983
rect 3598 939 3698 983
rect 144 513 244 573
rect 368 513 468 573
rect 582 513 682 573
rect 806 513 906 573
rect 144 500 906 513
rect 144 454 273 500
rect 319 454 497 500
rect 543 454 721 500
rect 767 454 906 500
rect 144 441 906 454
rect 144 377 244 441
rect 124 333 244 377
rect 348 333 468 441
rect 572 333 692 441
rect 796 377 906 441
rect 1030 500 1130 573
rect 1030 454 1071 500
rect 1117 454 1130 500
rect 1030 377 1130 454
rect 1254 513 1354 573
rect 1478 513 1578 573
rect 1712 513 1812 573
rect 1926 513 2026 573
rect 1254 500 1588 513
rect 1254 454 1529 500
rect 1575 454 1588 500
rect 1254 441 1588 454
rect 1254 377 1364 441
rect 796 333 916 377
rect 1020 333 1140 377
rect 1244 333 1364 377
rect 1468 333 1588 441
rect 1712 500 2026 513
rect 1712 454 1929 500
rect 1975 454 2026 500
rect 1712 441 2026 454
rect 1712 377 1812 441
rect 1692 333 1812 377
rect 1916 377 2026 441
rect 2150 513 2250 573
rect 2374 513 2474 573
rect 2150 500 2474 513
rect 2150 454 2163 500
rect 2209 454 2474 500
rect 2150 441 2474 454
rect 2150 377 2260 441
rect 1916 333 2036 377
rect 2140 333 2260 377
rect 2364 377 2474 441
rect 2588 500 2688 573
rect 2588 454 2601 500
rect 2647 454 2688 500
rect 2588 377 2688 454
rect 2936 513 3036 610
rect 3170 513 3270 610
rect 3374 513 3474 610
rect 3598 513 3698 610
rect 2936 500 3698 513
rect 2936 454 3065 500
rect 3111 454 3289 500
rect 3335 454 3513 500
rect 3559 454 3698 500
rect 2936 441 3698 454
rect 2936 377 3036 441
rect 2364 333 2484 377
rect 2588 333 2708 377
rect 2916 333 3036 377
rect 3140 333 3260 441
rect 3364 333 3484 441
rect 3588 377 3698 441
rect 3588 333 3708 377
rect 124 25 244 69
rect 348 25 468 69
rect 572 25 692 69
rect 796 25 916 69
rect 1020 25 1140 69
rect 1244 25 1364 69
rect 1468 25 1588 69
rect 1692 25 1812 69
rect 1916 25 2036 69
rect 2140 25 2260 69
rect 2364 25 2484 69
rect 2588 25 2708 69
rect 2916 25 3036 69
rect 3140 25 3260 69
rect 3364 25 3484 69
rect 3588 25 3708 69
<< polycontact >>
rect 273 454 319 500
rect 497 454 543 500
rect 721 454 767 500
rect 1071 454 1117 500
rect 1529 454 1575 500
rect 1929 454 1975 500
rect 2163 454 2209 500
rect 2601 454 2647 500
rect 3065 454 3111 500
rect 3289 454 3335 500
rect 3513 454 3559 500
<< metal1 >>
rect 0 926 3920 1098
rect 0 918 2861 926
rect 69 861 115 872
rect 69 664 115 721
rect 273 861 319 918
rect 273 710 319 721
rect 497 861 543 872
rect 497 664 543 721
rect 711 861 757 918
rect 711 710 757 721
rect 987 824 1841 870
rect 1887 824 2717 870
rect 2763 824 2774 870
rect 987 664 1033 824
rect 2907 918 3920 926
rect 1392 767 2325 778
rect 2861 775 2907 786
rect 3065 861 3111 872
rect 1392 721 1403 767
rect 1449 721 2279 767
rect 69 618 1033 664
rect 2279 684 2325 721
rect 3065 684 3111 721
rect 3299 861 3345 918
rect 3299 710 3345 721
rect 3503 861 3549 872
rect 2279 664 3111 684
rect 3503 664 3549 721
rect 3727 861 3773 918
rect 3727 710 3773 721
rect 2279 638 3549 664
rect 2693 618 3549 638
rect 1071 546 2647 592
rect 1071 500 1117 546
rect 1918 500 1986 546
rect 2601 500 2647 546
rect 254 454 273 500
rect 319 454 497 500
rect 543 454 721 500
rect 767 454 778 500
rect 1518 454 1529 500
rect 1575 454 1650 500
rect 1918 454 1929 500
rect 1975 454 1986 500
rect 2032 454 2163 500
rect 2209 454 2220 500
rect 254 354 306 454
rect 1071 443 1117 454
rect 1598 400 1650 454
rect 2032 400 2078 454
rect 2601 443 2647 454
rect 1598 354 2078 400
rect 2693 397 2739 618
rect 3054 500 3570 542
rect 3054 454 3065 500
rect 3111 454 3289 500
rect 3335 454 3513 500
rect 3559 454 3570 500
rect 2124 351 2739 397
rect 2785 362 3783 408
rect 49 312 95 323
rect 339 308 1565 321
rect 2124 308 2170 351
rect 273 285 2170 308
rect 319 275 2170 285
rect 319 239 372 275
rect 273 228 372 239
rect 710 274 778 275
rect 497 218 543 229
rect 710 228 721 274
rect 767 228 778 274
rect 1038 274 1226 275
rect 95 172 497 182
rect 945 218 991 229
rect 1038 228 1169 274
rect 1215 228 1226 274
rect 1532 274 2170 275
rect 543 172 945 182
rect 1393 218 1439 229
rect 1532 228 1617 274
rect 1663 262 2065 274
rect 1663 228 1674 262
rect 2054 228 2065 262
rect 2111 228 2170 274
rect 2289 294 2335 305
rect 991 172 1393 182
rect 1830 182 1841 216
rect 1439 172 1841 182
rect 49 170 1841 172
rect 1887 182 1898 216
rect 1887 170 2289 182
rect 49 154 2289 170
rect 2513 285 2559 351
rect 2513 228 2559 239
rect 2785 312 2831 362
rect 2335 172 2785 182
rect 2335 154 2831 172
rect 49 136 2831 154
rect 3065 305 3111 316
rect 3065 90 3111 165
rect 3289 312 3335 362
rect 3289 161 3335 172
rect 3513 305 3559 316
rect 3513 90 3559 165
rect 3737 312 3783 362
rect 3737 161 3783 172
rect 0 -90 3920 90
<< labels >>
flabel metal1 s 2032 454 2220 500 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 1071 546 2647 592 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 254 454 778 500 0 FreeSans 200 0 0 0 A3
port 3 nsew default input
flabel metal1 s 3054 454 3570 542 0 FreeSans 200 0 0 0 B
port 4 nsew default input
flabel metal1 s 0 918 3920 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 3513 90 3559 316 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 3503 778 3549 872 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 1518 454 1650 500 1 A1
port 1 nsew default input
rlabel metal1 s 2032 400 2078 454 1 A1
port 1 nsew default input
rlabel metal1 s 1598 400 1650 454 1 A1
port 1 nsew default input
rlabel metal1 s 1598 354 2078 400 1 A1
port 1 nsew default input
rlabel metal1 s 2601 454 2647 546 1 A2
port 2 nsew default input
rlabel metal1 s 1918 454 1986 546 1 A2
port 2 nsew default input
rlabel metal1 s 1071 454 1117 546 1 A2
port 2 nsew default input
rlabel metal1 s 2601 443 2647 454 1 A2
port 2 nsew default input
rlabel metal1 s 1071 443 1117 454 1 A2
port 2 nsew default input
rlabel metal1 s 254 354 306 454 1 A3
port 3 nsew default input
rlabel metal1 s 3065 778 3111 872 1 ZN
port 5 nsew default output
rlabel metal1 s 3503 721 3549 778 1 ZN
port 5 nsew default output
rlabel metal1 s 3065 721 3111 778 1 ZN
port 5 nsew default output
rlabel metal1 s 1392 721 2325 778 1 ZN
port 5 nsew default output
rlabel metal1 s 3503 684 3549 721 1 ZN
port 5 nsew default output
rlabel metal1 s 3065 684 3111 721 1 ZN
port 5 nsew default output
rlabel metal1 s 2279 684 2325 721 1 ZN
port 5 nsew default output
rlabel metal1 s 3503 664 3549 684 1 ZN
port 5 nsew default output
rlabel metal1 s 2279 664 3111 684 1 ZN
port 5 nsew default output
rlabel metal1 s 2279 638 3549 664 1 ZN
port 5 nsew default output
rlabel metal1 s 2693 618 3549 638 1 ZN
port 5 nsew default output
rlabel metal1 s 2693 397 2739 618 1 ZN
port 5 nsew default output
rlabel metal1 s 2124 351 2739 397 1 ZN
port 5 nsew default output
rlabel metal1 s 2513 321 2559 351 1 ZN
port 5 nsew default output
rlabel metal1 s 2124 321 2170 351 1 ZN
port 5 nsew default output
rlabel metal1 s 2513 308 2559 321 1 ZN
port 5 nsew default output
rlabel metal1 s 2124 308 2170 321 1 ZN
port 5 nsew default output
rlabel metal1 s 339 308 1565 321 1 ZN
port 5 nsew default output
rlabel metal1 s 2513 275 2559 308 1 ZN
port 5 nsew default output
rlabel metal1 s 273 275 2170 308 1 ZN
port 5 nsew default output
rlabel metal1 s 2513 262 2559 275 1 ZN
port 5 nsew default output
rlabel metal1 s 1532 262 2170 275 1 ZN
port 5 nsew default output
rlabel metal1 s 1038 262 1226 275 1 ZN
port 5 nsew default output
rlabel metal1 s 710 262 778 275 1 ZN
port 5 nsew default output
rlabel metal1 s 273 262 372 275 1 ZN
port 5 nsew default output
rlabel metal1 s 2513 228 2559 262 1 ZN
port 5 nsew default output
rlabel metal1 s 2054 228 2170 262 1 ZN
port 5 nsew default output
rlabel metal1 s 1532 228 1674 262 1 ZN
port 5 nsew default output
rlabel metal1 s 1038 228 1226 262 1 ZN
port 5 nsew default output
rlabel metal1 s 710 228 778 262 1 ZN
port 5 nsew default output
rlabel metal1 s 273 228 372 262 1 ZN
port 5 nsew default output
rlabel metal1 s 3727 775 3773 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3299 775 3345 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2861 775 2907 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 711 775 757 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 775 319 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3727 710 3773 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3299 710 3345 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 711 710 757 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 273 710 319 775 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3065 90 3111 316 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3920 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3920 1008
string GDS_END 158050
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 150130
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
