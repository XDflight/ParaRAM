magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -89 48 11 2153
rect 191 266 291 2153
rect 511 503 611 2153
rect 791 784 891 2153
rect 791 684 942 784
rect 511 403 717 503
rect 191 166 515 266
rect -89 -52 96 48
rect -4 -63 96 -52
rect 415 -63 515 166
rect 617 -63 717 403
rect 842 246 942 684
rect 1111 471 1211 2153
rect 1391 1010 1491 2153
rect 1391 910 1560 1010
rect 1111 371 1335 471
rect 842 146 1133 246
rect 1033 -63 1133 146
rect 1235 -63 1335 371
rect 1460 354 1560 910
rect 1711 630 1811 2153
rect 1991 858 2091 2153
rect 1991 758 2179 858
rect 1711 530 1955 630
rect 1460 254 1753 354
rect 1653 -63 1753 254
rect 1855 -63 1955 530
rect 2079 199 2179 758
rect 2311 404 2411 2153
rect 2591 619 2691 2153
rect 2911 821 3011 2153
rect 3191 1022 3291 2153
rect 3191 922 3360 1022
rect 2911 721 3193 821
rect 2591 519 2991 619
rect 2311 304 2574 404
rect 2079 99 2372 199
rect 2272 -63 2372 99
rect 2474 -63 2574 304
rect 2891 -63 2991 519
rect 3093 -63 3193 721
rect 3260 354 3360 922
rect 3511 565 3611 2153
rect 3791 850 3891 2153
rect 3791 750 4036 850
rect 3511 465 3813 565
rect 3260 254 3611 354
rect 3511 -63 3611 254
rect 3713 -63 3813 465
rect 3936 160 4036 750
rect 4111 320 4211 2153
rect 4391 847 4491 2153
rect 4391 747 4627 847
rect 4111 220 4431 320
rect 3936 60 4230 160
rect 4130 -63 4230 60
rect 4331 -63 4431 220
rect 4527 160 4627 747
rect 4527 60 4849 160
rect 4749 -63 4849 60
<< properties >>
string GDS_END 471110
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 469890
string path 13.205 10.765 13.205 2.845 14.705 2.845 14.705 -0.315 
<< end >>
