magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 4118 1094
<< pwell >>
rect -86 -86 4118 453
<< mvnmos >>
rect 248 69 368 306
rect 442 69 562 306
rect 666 69 786 306
rect 850 69 970 306
rect 1074 69 1194 306
rect 1258 69 1378 306
rect 1482 69 1602 306
rect 1666 69 1786 306
rect 1932 137 2052 295
rect 2156 137 2276 295
rect 2464 137 2584 295
rect 2688 137 2808 295
rect 2996 137 3116 295
rect 3220 137 3340 295
rect 3528 137 3648 295
rect 3752 137 3872 295
<< mvpmos >>
rect 258 573 358 939
rect 462 573 562 939
rect 666 573 766 939
rect 870 573 970 939
rect 1074 573 1174 939
rect 1278 573 1378 939
rect 1482 573 1582 939
rect 1686 573 1786 939
rect 1942 573 2042 939
rect 2166 573 2266 939
rect 2474 573 2574 939
rect 2698 573 2798 939
rect 3006 573 3106 939
rect 3230 573 3330 939
rect 3538 573 3638 939
rect 3762 573 3862 939
<< mvndiff >>
rect 122 222 248 306
rect 122 82 135 222
rect 181 82 248 222
rect 122 69 248 82
rect 368 69 442 306
rect 562 287 666 306
rect 562 147 591 287
rect 637 147 666 287
rect 562 69 666 147
rect 786 69 850 306
rect 970 128 1074 306
rect 970 82 999 128
rect 1045 82 1074 128
rect 970 69 1074 82
rect 1194 69 1258 306
rect 1378 293 1482 306
rect 1378 247 1407 293
rect 1453 247 1482 293
rect 1378 69 1482 247
rect 1602 69 1666 306
rect 1786 295 1866 306
rect 1786 190 1932 295
rect 1786 144 1815 190
rect 1861 144 1932 190
rect 1786 137 1932 144
rect 2052 282 2156 295
rect 2052 236 2081 282
rect 2127 236 2156 282
rect 2052 137 2156 236
rect 2276 190 2464 295
rect 2276 144 2347 190
rect 2393 144 2464 190
rect 2276 137 2464 144
rect 2584 282 2688 295
rect 2584 236 2613 282
rect 2659 236 2688 282
rect 2584 137 2688 236
rect 2808 190 2996 295
rect 2808 144 2879 190
rect 2925 144 2996 190
rect 2808 137 2996 144
rect 3116 282 3220 295
rect 3116 236 3145 282
rect 3191 236 3220 282
rect 3116 137 3220 236
rect 3340 190 3528 295
rect 3340 144 3411 190
rect 3457 144 3528 190
rect 3340 137 3528 144
rect 3648 282 3752 295
rect 3648 236 3677 282
rect 3723 236 3752 282
rect 3648 137 3752 236
rect 3872 196 3960 295
rect 3872 150 3901 196
rect 3947 150 3960 196
rect 3872 137 3960 150
rect 1786 69 1872 137
rect 2336 131 2404 137
rect 2868 131 2936 137
rect 3400 131 3468 137
<< mvpdiff >>
rect 170 861 258 939
rect 170 721 183 861
rect 229 721 258 861
rect 170 573 258 721
rect 358 769 462 939
rect 358 629 387 769
rect 433 629 462 769
rect 358 573 462 629
rect 562 861 666 939
rect 562 721 591 861
rect 637 721 666 861
rect 562 573 666 721
rect 766 769 870 939
rect 766 629 795 769
rect 841 629 870 769
rect 766 573 870 629
rect 970 861 1074 939
rect 970 721 999 861
rect 1045 721 1074 861
rect 970 573 1074 721
rect 1174 769 1278 939
rect 1174 629 1203 769
rect 1249 629 1278 769
rect 1174 573 1278 629
rect 1378 861 1482 939
rect 1378 721 1407 861
rect 1453 721 1482 861
rect 1378 573 1482 721
rect 1582 769 1686 939
rect 1582 629 1611 769
rect 1657 629 1686 769
rect 1582 573 1686 629
rect 1786 861 1942 939
rect 1786 721 1815 861
rect 1861 721 1942 861
rect 1786 573 1942 721
rect 2042 573 2166 939
rect 2266 881 2474 939
rect 2266 741 2295 881
rect 2341 741 2474 881
rect 2266 573 2474 741
rect 2574 573 2698 939
rect 2798 861 3006 939
rect 2798 721 2827 861
rect 2873 721 3006 861
rect 2798 573 3006 721
rect 3106 573 3230 939
rect 3330 881 3538 939
rect 3330 741 3359 881
rect 3405 741 3538 881
rect 3330 573 3538 741
rect 3638 573 3762 939
rect 3862 861 3950 939
rect 3862 721 3891 861
rect 3937 721 3950 861
rect 3862 573 3950 721
<< mvndiffc >>
rect 135 82 181 222
rect 591 147 637 287
rect 999 82 1045 128
rect 1407 247 1453 293
rect 1815 144 1861 190
rect 2081 236 2127 282
rect 2347 144 2393 190
rect 2613 236 2659 282
rect 2879 144 2925 190
rect 3145 236 3191 282
rect 3411 144 3457 190
rect 3677 236 3723 282
rect 3901 150 3947 196
<< mvpdiffc >>
rect 183 721 229 861
rect 387 629 433 769
rect 591 721 637 861
rect 795 629 841 769
rect 999 721 1045 861
rect 1203 629 1249 769
rect 1407 721 1453 861
rect 1611 629 1657 769
rect 1815 721 1861 861
rect 2295 741 2341 881
rect 2827 721 2873 861
rect 3359 741 3405 881
rect 3891 721 3937 861
<< polysilicon >>
rect 258 939 358 983
rect 462 939 562 983
rect 666 939 766 983
rect 870 939 970 983
rect 1074 939 1174 983
rect 1278 939 1378 983
rect 1482 939 1582 983
rect 1686 939 1786 983
rect 1942 939 2042 983
rect 2166 939 2266 983
rect 2474 939 2574 983
rect 2698 939 2798 983
rect 3006 939 3106 983
rect 3230 939 3330 983
rect 3538 939 3638 983
rect 3762 939 3862 983
rect 258 513 358 573
rect 462 513 562 573
rect 666 513 766 573
rect 258 500 368 513
rect 258 454 309 500
rect 355 454 368 500
rect 258 350 368 454
rect 462 491 766 513
rect 870 513 970 573
rect 1074 513 1174 573
rect 870 500 1174 513
rect 462 480 786 491
rect 462 441 713 480
rect 462 350 562 441
rect 248 306 368 350
rect 442 306 562 350
rect 666 434 713 441
rect 759 434 786 480
rect 666 306 786 434
rect 870 454 1023 500
rect 1069 454 1174 500
rect 1278 513 1378 573
rect 1482 513 1582 573
rect 1278 493 1582 513
rect 870 441 1174 454
rect 870 350 970 441
rect 850 306 970 350
rect 1074 350 1174 441
rect 1258 480 1582 493
rect 1258 434 1271 480
rect 1317 441 1582 480
rect 1317 434 1378 441
rect 1074 306 1194 350
rect 1258 306 1378 434
rect 1482 350 1582 441
rect 1686 500 1786 573
rect 1686 454 1699 500
rect 1745 454 1786 500
rect 1686 350 1786 454
rect 1482 306 1602 350
rect 1666 306 1786 350
rect 1942 500 2042 573
rect 1942 454 1983 500
rect 2029 454 2042 500
rect 1942 339 2042 454
rect 2166 513 2266 573
rect 2474 513 2574 573
rect 2698 513 2798 573
rect 3006 513 3106 573
rect 2166 500 2574 513
rect 2166 454 2515 500
rect 2561 454 2574 500
rect 2166 441 2574 454
rect 2166 339 2276 441
rect 1932 295 2052 339
rect 2156 295 2276 339
rect 2464 339 2574 441
rect 2688 500 3106 513
rect 2688 454 2701 500
rect 2747 454 3106 500
rect 2688 441 3106 454
rect 2464 295 2584 339
rect 2688 295 2808 441
rect 2996 339 3106 441
rect 3230 513 3330 573
rect 3538 513 3638 573
rect 3230 500 3638 513
rect 3230 454 3243 500
rect 3289 454 3638 500
rect 3230 441 3638 454
rect 3230 339 3340 441
rect 2996 295 3116 339
rect 3220 295 3340 339
rect 3528 339 3638 441
rect 3762 500 3862 573
rect 3762 454 3803 500
rect 3849 454 3862 500
rect 3762 339 3862 454
rect 3528 295 3648 339
rect 3752 295 3872 339
rect 1932 93 2052 137
rect 2156 93 2276 137
rect 2464 93 2584 137
rect 2688 93 2808 137
rect 2996 93 3116 137
rect 3220 93 3340 137
rect 3528 93 3648 137
rect 3752 93 3872 137
rect 248 25 368 69
rect 442 25 562 69
rect 666 25 786 69
rect 850 25 970 69
rect 1074 25 1194 69
rect 1258 25 1378 69
rect 1482 25 1602 69
rect 1666 25 1786 69
<< polycontact >>
rect 309 454 355 500
rect 713 434 759 480
rect 1023 454 1069 500
rect 1271 434 1317 480
rect 1699 454 1745 500
rect 1983 454 2029 500
rect 2515 454 2561 500
rect 2701 454 2747 500
rect 3243 454 3289 500
rect 3803 454 3849 500
<< metal1 >>
rect 0 918 4032 1098
rect 2295 881 2341 918
rect 183 861 1861 872
rect 229 826 591 861
rect 183 710 229 721
rect 387 769 433 780
rect 217 629 387 664
rect 637 826 999 861
rect 591 710 637 721
rect 795 769 841 780
rect 433 629 795 664
rect 1045 826 1407 861
rect 999 710 1045 721
rect 1150 769 1249 780
rect 1150 664 1203 769
rect 841 629 1203 664
rect 1453 826 1815 861
rect 1407 710 1453 721
rect 1611 769 1657 780
rect 1249 629 1611 664
rect 3359 881 3405 918
rect 2295 730 2341 741
rect 2827 861 2873 872
rect 1815 684 1861 721
rect 3359 730 3405 741
rect 3891 861 3937 872
rect 2827 684 2873 721
rect 3891 684 3937 721
rect 1815 638 3937 684
rect 217 618 1657 629
rect 217 308 263 618
rect 309 526 1745 572
rect 309 500 355 526
rect 1023 500 1069 526
rect 309 443 355 454
rect 702 434 713 480
rect 759 434 770 480
rect 1374 500 1745 526
rect 1023 443 1069 454
rect 702 430 770 434
rect 1115 434 1271 480
rect 1317 434 1328 480
rect 1374 454 1699 500
rect 1972 546 3890 592
rect 1972 500 2040 546
rect 2701 500 2747 546
rect 3792 500 3890 546
rect 1972 454 1983 500
rect 2029 454 2040 500
rect 2504 454 2515 500
rect 2561 454 2572 500
rect 1374 443 1745 454
rect 702 397 978 430
rect 1115 397 1161 434
rect 702 351 1161 397
rect 2504 397 2572 454
rect 2701 443 2747 454
rect 2838 454 3243 500
rect 3289 454 3300 500
rect 3792 454 3803 500
rect 3849 454 3890 500
rect 2838 430 2884 454
rect 2792 397 2884 430
rect 2504 351 2884 397
rect 217 305 608 308
rect 217 293 3734 305
rect 217 287 1407 293
rect 217 262 591 287
rect 135 222 181 233
rect 0 82 135 90
rect 637 247 1407 287
rect 1453 282 3734 293
rect 1453 247 2081 282
rect 637 236 2081 247
rect 2127 236 2613 282
rect 2659 236 3145 282
rect 3191 236 3677 282
rect 3723 236 3734 282
rect 3901 196 3947 207
rect 591 136 637 147
rect 1804 144 1815 190
rect 1861 144 1872 190
rect 999 128 1045 139
rect 181 82 999 90
rect 1804 90 1872 144
rect 2336 144 2347 190
rect 2393 144 2404 190
rect 2336 90 2404 144
rect 2868 144 2879 190
rect 2925 144 2936 190
rect 2868 90 2936 144
rect 3400 144 3411 190
rect 3457 144 3468 190
rect 3400 90 3468 144
rect 3901 90 3947 150
rect 1045 82 4032 90
rect 0 -90 4032 82
<< labels >>
flabel metal1 s 1115 434 1328 480 0 FreeSans 200 0 0 0 A1
port 1 nsew default input
flabel metal1 s 309 526 1745 572 0 FreeSans 200 0 0 0 A2
port 2 nsew default input
flabel metal1 s 1972 546 3890 592 0 FreeSans 200 0 0 0 B
port 3 nsew default input
flabel metal1 s 2838 454 3300 500 0 FreeSans 200 0 0 0 C
port 4 nsew default input
flabel metal1 s 0 918 4032 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 135 207 181 233 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel metal1 s 1611 664 1657 780 0 FreeSans 200 0 0 0 ZN
port 5 nsew default output
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 702 434 770 480 1 A1
port 1 nsew default input
rlabel metal1 s 1115 430 1161 434 1 A1
port 1 nsew default input
rlabel metal1 s 702 430 770 434 1 A1
port 1 nsew default input
rlabel metal1 s 1115 397 1161 430 1 A1
port 1 nsew default input
rlabel metal1 s 702 397 978 430 1 A1
port 1 nsew default input
rlabel metal1 s 702 351 1161 397 1 A1
port 1 nsew default input
rlabel metal1 s 1374 443 1745 526 1 A2
port 2 nsew default input
rlabel metal1 s 1023 443 1069 526 1 A2
port 2 nsew default input
rlabel metal1 s 309 443 355 526 1 A2
port 2 nsew default input
rlabel metal1 s 3792 454 3890 546 1 B
port 3 nsew default input
rlabel metal1 s 2701 454 2747 546 1 B
port 3 nsew default input
rlabel metal1 s 1972 454 2040 546 1 B
port 3 nsew default input
rlabel metal1 s 2701 443 2747 454 1 B
port 3 nsew default input
rlabel metal1 s 2504 454 2572 500 1 C
port 4 nsew default input
rlabel metal1 s 2838 430 2884 454 1 C
port 4 nsew default input
rlabel metal1 s 2504 430 2572 454 1 C
port 4 nsew default input
rlabel metal1 s 2792 397 2884 430 1 C
port 4 nsew default input
rlabel metal1 s 2504 397 2572 430 1 C
port 4 nsew default input
rlabel metal1 s 2504 351 2884 397 1 C
port 4 nsew default input
rlabel metal1 s 1150 664 1249 780 1 ZN
port 5 nsew default output
rlabel metal1 s 795 664 841 780 1 ZN
port 5 nsew default output
rlabel metal1 s 387 664 433 780 1 ZN
port 5 nsew default output
rlabel metal1 s 217 618 1657 664 1 ZN
port 5 nsew default output
rlabel metal1 s 217 308 263 618 1 ZN
port 5 nsew default output
rlabel metal1 s 217 305 608 308 1 ZN
port 5 nsew default output
rlabel metal1 s 217 262 3734 305 1 ZN
port 5 nsew default output
rlabel metal1 s 591 236 3734 262 1 ZN
port 5 nsew default output
rlabel metal1 s 591 136 637 236 1 ZN
port 5 nsew default output
rlabel metal1 s 3359 730 3405 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2295 730 2341 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3901 190 3947 207 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 135 190 181 207 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3901 139 3947 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3400 139 3468 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2868 139 2936 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2336 139 2404 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1804 139 1872 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 135 139 181 190 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3901 90 3947 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3400 90 3468 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2868 90 2936 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2336 90 2404 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1804 90 1872 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 999 90 1045 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 135 90 181 139 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4032 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 1008
string GDS_END 1191386
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1183882
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
