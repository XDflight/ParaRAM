magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 343 -141
<< polysilicon >>
rect -31 2631 88 2703
rect -31 -73 88 -1
use pmos_5p04310590878171_256x8m81  pmos_5p04310590878171_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 2752
<< properties >>
string GDS_END 292958
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 292644
<< end >>
