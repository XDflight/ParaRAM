magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -81 819 81 825
rect -81 793 -75 819
rect -49 793 -13 819
rect 13 793 49 819
rect 75 793 81 819
rect -81 757 81 793
rect -81 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 81 757
rect -81 695 81 731
rect -81 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 81 695
rect -81 633 81 669
rect -81 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 81 633
rect -81 571 81 607
rect -81 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 81 571
rect -81 509 81 545
rect -81 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 81 509
rect -81 447 81 483
rect -81 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 81 447
rect -81 385 81 421
rect -81 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 81 385
rect -81 323 81 359
rect -81 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 81 323
rect -81 261 81 297
rect -81 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 81 261
rect -81 199 81 235
rect -81 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 81 199
rect -81 137 81 173
rect -81 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 81 137
rect -81 75 81 111
rect -81 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 81 75
rect -81 13 81 49
rect -81 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 81 13
rect -81 -49 81 -13
rect -81 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 81 -49
rect -81 -111 81 -75
rect -81 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 81 -111
rect -81 -173 81 -137
rect -81 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 81 -173
rect -81 -235 81 -199
rect -81 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 81 -235
rect -81 -297 81 -261
rect -81 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 81 -297
rect -81 -359 81 -323
rect -81 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 81 -359
rect -81 -421 81 -385
rect -81 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 81 -421
rect -81 -483 81 -447
rect -81 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 81 -483
rect -81 -545 81 -509
rect -81 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 81 -545
rect -81 -607 81 -571
rect -81 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 81 -607
rect -81 -669 81 -633
rect -81 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 81 -669
rect -81 -731 81 -695
rect -81 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 81 -731
rect -81 -793 81 -757
rect -81 -819 -75 -793
rect -49 -819 -13 -793
rect 13 -819 49 -793
rect 75 -819 81 -793
rect -81 -825 81 -819
<< via1 >>
rect -75 793 -49 819
rect -13 793 13 819
rect 49 793 75 819
rect -75 731 -49 757
rect -13 731 13 757
rect 49 731 75 757
rect -75 669 -49 695
rect -13 669 13 695
rect 49 669 75 695
rect -75 607 -49 633
rect -13 607 13 633
rect 49 607 75 633
rect -75 545 -49 571
rect -13 545 13 571
rect 49 545 75 571
rect -75 483 -49 509
rect -13 483 13 509
rect 49 483 75 509
rect -75 421 -49 447
rect -13 421 13 447
rect 49 421 75 447
rect -75 359 -49 385
rect -13 359 13 385
rect 49 359 75 385
rect -75 297 -49 323
rect -13 297 13 323
rect 49 297 75 323
rect -75 235 -49 261
rect -13 235 13 261
rect 49 235 75 261
rect -75 173 -49 199
rect -13 173 13 199
rect 49 173 75 199
rect -75 111 -49 137
rect -13 111 13 137
rect 49 111 75 137
rect -75 49 -49 75
rect -13 49 13 75
rect 49 49 75 75
rect -75 -13 -49 13
rect -13 -13 13 13
rect 49 -13 75 13
rect -75 -75 -49 -49
rect -13 -75 13 -49
rect 49 -75 75 -49
rect -75 -137 -49 -111
rect -13 -137 13 -111
rect 49 -137 75 -111
rect -75 -199 -49 -173
rect -13 -199 13 -173
rect 49 -199 75 -173
rect -75 -261 -49 -235
rect -13 -261 13 -235
rect 49 -261 75 -235
rect -75 -323 -49 -297
rect -13 -323 13 -297
rect 49 -323 75 -297
rect -75 -385 -49 -359
rect -13 -385 13 -359
rect 49 -385 75 -359
rect -75 -447 -49 -421
rect -13 -447 13 -421
rect 49 -447 75 -421
rect -75 -509 -49 -483
rect -13 -509 13 -483
rect 49 -509 75 -483
rect -75 -571 -49 -545
rect -13 -571 13 -545
rect 49 -571 75 -545
rect -75 -633 -49 -607
rect -13 -633 13 -607
rect 49 -633 75 -607
rect -75 -695 -49 -669
rect -13 -695 13 -669
rect 49 -695 75 -669
rect -75 -757 -49 -731
rect -13 -757 13 -731
rect 49 -757 75 -731
rect -75 -819 -49 -793
rect -13 -819 13 -793
rect 49 -819 75 -793
<< metal2 >>
rect -81 819 81 825
rect -81 793 -75 819
rect -49 793 -13 819
rect 13 793 49 819
rect 75 793 81 819
rect -81 757 81 793
rect -81 731 -75 757
rect -49 731 -13 757
rect 13 731 49 757
rect 75 731 81 757
rect -81 695 81 731
rect -81 669 -75 695
rect -49 669 -13 695
rect 13 669 49 695
rect 75 669 81 695
rect -81 633 81 669
rect -81 607 -75 633
rect -49 607 -13 633
rect 13 607 49 633
rect 75 607 81 633
rect -81 571 81 607
rect -81 545 -75 571
rect -49 545 -13 571
rect 13 545 49 571
rect 75 545 81 571
rect -81 509 81 545
rect -81 483 -75 509
rect -49 483 -13 509
rect 13 483 49 509
rect 75 483 81 509
rect -81 447 81 483
rect -81 421 -75 447
rect -49 421 -13 447
rect 13 421 49 447
rect 75 421 81 447
rect -81 385 81 421
rect -81 359 -75 385
rect -49 359 -13 385
rect 13 359 49 385
rect 75 359 81 385
rect -81 323 81 359
rect -81 297 -75 323
rect -49 297 -13 323
rect 13 297 49 323
rect 75 297 81 323
rect -81 261 81 297
rect -81 235 -75 261
rect -49 235 -13 261
rect 13 235 49 261
rect 75 235 81 261
rect -81 199 81 235
rect -81 173 -75 199
rect -49 173 -13 199
rect 13 173 49 199
rect 75 173 81 199
rect -81 137 81 173
rect -81 111 -75 137
rect -49 111 -13 137
rect 13 111 49 137
rect 75 111 81 137
rect -81 75 81 111
rect -81 49 -75 75
rect -49 49 -13 75
rect 13 49 49 75
rect 75 49 81 75
rect -81 13 81 49
rect -81 -13 -75 13
rect -49 -13 -13 13
rect 13 -13 49 13
rect 75 -13 81 13
rect -81 -49 81 -13
rect -81 -75 -75 -49
rect -49 -75 -13 -49
rect 13 -75 49 -49
rect 75 -75 81 -49
rect -81 -111 81 -75
rect -81 -137 -75 -111
rect -49 -137 -13 -111
rect 13 -137 49 -111
rect 75 -137 81 -111
rect -81 -173 81 -137
rect -81 -199 -75 -173
rect -49 -199 -13 -173
rect 13 -199 49 -173
rect 75 -199 81 -173
rect -81 -235 81 -199
rect -81 -261 -75 -235
rect -49 -261 -13 -235
rect 13 -261 49 -235
rect 75 -261 81 -235
rect -81 -297 81 -261
rect -81 -323 -75 -297
rect -49 -323 -13 -297
rect 13 -323 49 -297
rect 75 -323 81 -297
rect -81 -359 81 -323
rect -81 -385 -75 -359
rect -49 -385 -13 -359
rect 13 -385 49 -359
rect 75 -385 81 -359
rect -81 -421 81 -385
rect -81 -447 -75 -421
rect -49 -447 -13 -421
rect 13 -447 49 -421
rect 75 -447 81 -421
rect -81 -483 81 -447
rect -81 -509 -75 -483
rect -49 -509 -13 -483
rect 13 -509 49 -483
rect 75 -509 81 -483
rect -81 -545 81 -509
rect -81 -571 -75 -545
rect -49 -571 -13 -545
rect 13 -571 49 -545
rect 75 -571 81 -545
rect -81 -607 81 -571
rect -81 -633 -75 -607
rect -49 -633 -13 -607
rect 13 -633 49 -607
rect 75 -633 81 -607
rect -81 -669 81 -633
rect -81 -695 -75 -669
rect -49 -695 -13 -669
rect 13 -695 49 -669
rect 75 -695 81 -669
rect -81 -731 81 -695
rect -81 -757 -75 -731
rect -49 -757 -13 -731
rect 13 -757 49 -731
rect 75 -757 81 -731
rect -81 -793 81 -757
rect -81 -819 -75 -793
rect -49 -819 -13 -793
rect 13 -819 49 -793
rect 75 -819 81 -793
rect -81 -825 81 -819
<< properties >>
string GDS_END 733312
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 727996
<< end >>
