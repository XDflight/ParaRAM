magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -2038 -390 2039 391
<< nsubdiff >>
rect -1895 186 1896 244
rect -1895 140 -1841 186
rect -1795 140 -1683 186
rect -1637 140 -1525 186
rect -1479 140 -1367 186
rect -1321 140 -1209 186
rect -1163 140 -1051 186
rect -1005 140 -893 186
rect -847 140 -735 186
rect -689 140 -577 186
rect -531 140 -418 186
rect -372 140 -260 186
rect -214 140 -102 186
rect -56 140 56 186
rect 102 140 214 186
rect 260 140 372 186
rect 418 140 531 186
rect 577 140 689 186
rect 735 140 847 186
rect 893 140 1005 186
rect 1051 140 1163 186
rect 1209 140 1321 186
rect 1367 140 1479 186
rect 1525 140 1637 186
rect 1683 140 1795 186
rect 1841 140 1896 186
rect -1895 23 1896 140
rect -1895 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1896 23
rect -1895 -140 1896 -23
rect -1895 -186 -1841 -140
rect -1795 -186 -1683 -140
rect -1637 -186 -1525 -140
rect -1479 -186 -1367 -140
rect -1321 -186 -1209 -140
rect -1163 -186 -1051 -140
rect -1005 -186 -893 -140
rect -847 -186 -735 -140
rect -689 -186 -577 -140
rect -531 -186 -418 -140
rect -372 -186 -260 -140
rect -214 -186 -102 -140
rect -56 -186 56 -140
rect 102 -186 214 -140
rect 260 -186 372 -140
rect 418 -186 531 -140
rect 577 -186 689 -140
rect 735 -186 847 -140
rect 893 -186 1005 -140
rect 1051 -186 1163 -140
rect 1209 -186 1321 -140
rect 1367 -186 1479 -140
rect 1525 -186 1637 -140
rect 1683 -186 1795 -140
rect 1841 -186 1896 -140
rect -1895 -243 1896 -186
<< nsubdiffcont >>
rect -1841 140 -1795 186
rect -1683 140 -1637 186
rect -1525 140 -1479 186
rect -1367 140 -1321 186
rect -1209 140 -1163 186
rect -1051 140 -1005 186
rect -893 140 -847 186
rect -735 140 -689 186
rect -577 140 -531 186
rect -418 140 -372 186
rect -260 140 -214 186
rect -102 140 -56 186
rect 56 140 102 186
rect 214 140 260 186
rect 372 140 418 186
rect 531 140 577 186
rect 689 140 735 186
rect 847 140 893 186
rect 1005 140 1051 186
rect 1163 140 1209 186
rect 1321 140 1367 186
rect 1479 140 1525 186
rect 1637 140 1683 186
rect 1795 140 1841 186
rect -1841 -23 -1795 23
rect -1683 -23 -1637 23
rect -1525 -23 -1479 23
rect -1367 -23 -1321 23
rect -1209 -23 -1163 23
rect -1051 -23 -1005 23
rect -893 -23 -847 23
rect -735 -23 -689 23
rect -577 -23 -531 23
rect -418 -23 -372 23
rect -260 -23 -214 23
rect -102 -23 -56 23
rect 56 -23 102 23
rect 214 -23 260 23
rect 372 -23 418 23
rect 531 -23 577 23
rect 689 -23 735 23
rect 847 -23 893 23
rect 1005 -23 1051 23
rect 1163 -23 1209 23
rect 1321 -23 1367 23
rect 1479 -23 1525 23
rect 1637 -23 1683 23
rect 1795 -23 1841 23
rect -1841 -186 -1795 -140
rect -1683 -186 -1637 -140
rect -1525 -186 -1479 -140
rect -1367 -186 -1321 -140
rect -1209 -186 -1163 -140
rect -1051 -186 -1005 -140
rect -893 -186 -847 -140
rect -735 -186 -689 -140
rect -577 -186 -531 -140
rect -418 -186 -372 -140
rect -260 -186 -214 -140
rect -102 -186 -56 -140
rect 56 -186 102 -140
rect 214 -186 260 -140
rect 372 -186 418 -140
rect 531 -186 577 -140
rect 689 -186 735 -140
rect 847 -186 893 -140
rect 1005 -186 1051 -140
rect 1163 -186 1209 -140
rect 1321 -186 1367 -140
rect 1479 -186 1525 -140
rect 1637 -186 1683 -140
rect 1795 -186 1841 -140
<< metal1 >>
rect -1876 186 1876 223
rect -1876 140 -1841 186
rect -1795 140 -1683 186
rect -1637 140 -1525 186
rect -1479 140 -1367 186
rect -1321 140 -1209 186
rect -1163 140 -1051 186
rect -1005 140 -893 186
rect -847 140 -735 186
rect -689 140 -577 186
rect -531 140 -418 186
rect -372 140 -260 186
rect -214 140 -102 186
rect -56 140 56 186
rect 102 140 214 186
rect 260 140 372 186
rect 418 140 531 186
rect 577 140 689 186
rect 735 140 847 186
rect 893 140 1005 186
rect 1051 140 1163 186
rect 1209 140 1321 186
rect 1367 140 1479 186
rect 1525 140 1637 186
rect 1683 140 1795 186
rect 1841 140 1876 186
rect -1876 23 1876 140
rect -1876 -23 -1841 23
rect -1795 -23 -1683 23
rect -1637 -23 -1525 23
rect -1479 -23 -1367 23
rect -1321 -23 -1209 23
rect -1163 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1163 23
rect 1209 -23 1321 23
rect 1367 -23 1479 23
rect 1525 -23 1637 23
rect 1683 -23 1795 23
rect 1841 -23 1876 23
rect -1876 -140 1876 -23
rect -1876 -186 -1841 -140
rect -1795 -186 -1683 -140
rect -1637 -186 -1525 -140
rect -1479 -186 -1367 -140
rect -1321 -186 -1209 -140
rect -1163 -186 -1051 -140
rect -1005 -186 -893 -140
rect -847 -186 -735 -140
rect -689 -186 -577 -140
rect -531 -186 -418 -140
rect -372 -186 -260 -140
rect -214 -186 -102 -140
rect -56 -186 56 -140
rect 102 -186 214 -140
rect 260 -186 372 -140
rect 418 -186 531 -140
rect 577 -186 689 -140
rect 735 -186 847 -140
rect 893 -186 1005 -140
rect 1051 -186 1163 -140
rect 1209 -186 1321 -140
rect 1367 -186 1479 -140
rect 1525 -186 1637 -140
rect 1683 -186 1795 -140
rect 1841 -186 1876 -140
rect -1876 -223 1876 -186
<< properties >>
string GDS_END 650942
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 646074
<< end >>
