magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 3894 1094
<< pwell >>
rect -86 -86 3894 453
<< mvnmos >>
rect 132 69 252 333
rect 356 69 476 333
rect 624 173 744 333
rect 792 173 912 333
rect 960 173 1080 333
rect 1184 173 1304 333
rect 1408 173 1528 333
rect 1632 173 1752 333
rect 1856 173 1976 333
rect 2224 173 2344 333
rect 2448 173 2568 333
rect 2672 173 2792 333
rect 2896 173 3016 333
rect 3064 173 3184 333
rect 3328 69 3448 333
rect 3552 69 3672 333
<< mvpmos >>
rect 196 573 296 933
rect 400 573 500 933
rect 664 573 764 851
rect 812 573 912 851
rect 980 573 1080 851
rect 1184 573 1284 851
rect 1428 573 1528 851
rect 1632 573 1732 851
rect 1876 573 1976 851
rect 2224 573 2324 851
rect 2448 573 2548 851
rect 2692 573 2792 851
rect 2916 573 3016 851
rect 3064 573 3164 851
rect 3304 573 3404 933
rect 3508 573 3608 933
<< mvndiff >>
rect 44 222 132 333
rect 44 82 57 222
rect 103 82 132 222
rect 44 69 132 82
rect 252 320 356 333
rect 252 180 281 320
rect 327 180 356 320
rect 252 69 356 180
rect 476 222 624 333
rect 476 82 505 222
rect 551 173 624 222
rect 744 173 792 333
rect 912 173 960 333
rect 1080 320 1184 333
rect 1080 274 1109 320
rect 1155 274 1184 320
rect 1080 173 1184 274
rect 1304 320 1408 333
rect 1304 274 1333 320
rect 1379 274 1408 320
rect 1304 173 1408 274
rect 1528 232 1632 333
rect 1528 186 1557 232
rect 1603 186 1632 232
rect 1528 173 1632 186
rect 1752 320 1856 333
rect 1752 274 1781 320
rect 1827 274 1856 320
rect 1752 173 1856 274
rect 1976 232 2064 333
rect 1976 186 2005 232
rect 2051 186 2064 232
rect 1976 173 2064 186
rect 2136 320 2224 333
rect 2136 274 2149 320
rect 2195 274 2224 320
rect 2136 173 2224 274
rect 2344 232 2448 333
rect 2344 186 2373 232
rect 2419 186 2448 232
rect 2344 173 2448 186
rect 2568 320 2672 333
rect 2568 274 2597 320
rect 2643 274 2672 320
rect 2568 173 2672 274
rect 2792 320 2896 333
rect 2792 274 2821 320
rect 2867 274 2896 320
rect 2792 173 2896 274
rect 3016 173 3064 333
rect 3184 228 3328 333
rect 3184 182 3253 228
rect 3299 182 3328 228
rect 3184 173 3328 182
rect 551 82 564 173
rect 476 69 564 82
rect 3244 69 3328 173
rect 3448 320 3552 333
rect 3448 180 3477 320
rect 3523 180 3552 320
rect 3448 69 3552 180
rect 3672 222 3760 333
rect 3672 82 3701 222
rect 3747 82 3760 222
rect 3672 69 3760 82
<< mvpdiff >>
rect 108 920 196 933
rect 108 780 121 920
rect 167 780 196 920
rect 108 573 196 780
rect 296 726 400 933
rect 296 586 325 726
rect 371 586 400 726
rect 296 573 400 586
rect 500 920 588 933
rect 500 780 529 920
rect 575 851 588 920
rect 3224 851 3304 933
rect 575 780 664 851
rect 500 573 664 780
rect 764 573 812 851
rect 912 573 980 851
rect 1080 726 1184 851
rect 1080 586 1109 726
rect 1155 586 1184 726
rect 1080 573 1184 586
rect 1284 632 1428 851
rect 1284 586 1353 632
rect 1399 586 1428 632
rect 1284 573 1428 586
rect 1528 838 1632 851
rect 1528 792 1557 838
rect 1603 792 1632 838
rect 1528 573 1632 792
rect 1732 737 1876 851
rect 1732 597 1761 737
rect 1807 597 1876 737
rect 1732 573 1876 597
rect 1976 838 2064 851
rect 1976 698 2005 838
rect 2051 698 2064 838
rect 1976 573 2064 698
rect 2136 737 2224 851
rect 2136 597 2149 737
rect 2195 597 2224 737
rect 2136 573 2224 597
rect 2324 838 2448 851
rect 2324 698 2353 838
rect 2399 698 2448 838
rect 2324 573 2448 698
rect 2548 737 2692 851
rect 2548 597 2577 737
rect 2623 597 2692 737
rect 2548 573 2692 597
rect 2792 632 2916 851
rect 2792 586 2821 632
rect 2867 586 2916 632
rect 2792 573 2916 586
rect 3016 573 3064 851
rect 3164 838 3304 851
rect 3164 792 3193 838
rect 3239 792 3304 838
rect 3164 573 3304 792
rect 3404 726 3508 933
rect 3404 586 3433 726
rect 3479 586 3508 726
rect 3404 573 3508 586
rect 3608 920 3696 933
rect 3608 780 3637 920
rect 3683 780 3696 920
rect 3608 573 3696 780
<< mvndiffc >>
rect 57 82 103 222
rect 281 180 327 320
rect 505 82 551 222
rect 1109 274 1155 320
rect 1333 274 1379 320
rect 1557 186 1603 232
rect 1781 274 1827 320
rect 2005 186 2051 232
rect 2149 274 2195 320
rect 2373 186 2419 232
rect 2597 274 2643 320
rect 2821 274 2867 320
rect 3253 182 3299 228
rect 3477 180 3523 320
rect 3701 82 3747 222
<< mvpdiffc >>
rect 121 780 167 920
rect 325 586 371 726
rect 529 780 575 920
rect 1109 586 1155 726
rect 1353 586 1399 632
rect 1557 792 1603 838
rect 1761 597 1807 737
rect 2005 698 2051 838
rect 2149 597 2195 737
rect 2353 698 2399 838
rect 2577 597 2623 737
rect 2821 586 2867 632
rect 3193 792 3239 838
rect 3433 586 3479 726
rect 3637 780 3683 920
<< polysilicon >>
rect 196 933 296 977
rect 400 933 500 977
rect 812 943 3016 983
rect 664 851 764 895
rect 812 851 912 943
rect 980 851 1080 895
rect 1184 851 1284 895
rect 1428 851 1528 895
rect 1632 851 1732 943
rect 1876 851 1976 895
rect 2224 851 2324 943
rect 2448 851 2548 895
rect 2692 851 2792 895
rect 2916 851 3016 943
rect 3304 933 3404 977
rect 3508 933 3608 977
rect 3064 851 3164 895
rect 196 513 296 573
rect 400 529 500 573
rect 664 529 764 573
rect 400 513 476 529
rect 196 441 476 513
rect 196 377 252 441
rect 132 333 252 377
rect 356 412 476 441
rect 356 366 417 412
rect 463 366 476 412
rect 664 523 744 529
rect 664 477 685 523
rect 731 477 744 523
rect 664 377 744 477
rect 812 377 912 573
rect 980 430 1080 573
rect 980 384 1021 430
rect 1067 384 1080 430
rect 980 377 1080 384
rect 356 333 476 366
rect 624 333 744 377
rect 792 333 912 377
rect 960 333 1080 377
rect 1184 540 1284 573
rect 1184 494 1225 540
rect 1271 494 1284 540
rect 1184 377 1284 494
rect 1428 377 1528 573
rect 1184 333 1304 377
rect 1408 333 1528 377
rect 1632 377 1732 573
rect 1876 430 1976 573
rect 1876 384 1889 430
rect 1935 384 1976 430
rect 1876 377 1976 384
rect 1632 333 1752 377
rect 1856 333 1976 377
rect 2224 377 2324 573
rect 2448 377 2548 573
rect 2692 412 2792 573
rect 2692 377 2724 412
rect 2224 333 2344 377
rect 2448 333 2568 377
rect 2672 366 2724 377
rect 2770 366 2792 412
rect 2916 487 3016 573
rect 2916 441 2942 487
rect 2988 441 3016 487
rect 2916 377 3016 441
rect 2672 333 2792 366
rect 2896 333 3016 377
rect 3064 377 3164 573
rect 3304 513 3404 573
rect 3508 513 3608 573
rect 3328 508 3608 513
rect 3064 333 3184 377
rect 3328 366 3341 508
rect 3387 441 3608 508
rect 3387 366 3448 441
rect 3328 333 3448 366
rect 3552 377 3608 441
rect 3552 333 3672 377
rect 624 81 744 173
rect 792 129 912 173
rect 960 129 1080 173
rect 1184 129 1304 173
rect 1408 81 1528 173
rect 1632 129 1752 173
rect 1856 129 1976 173
rect 2224 129 2344 173
rect 2448 81 2568 173
rect 2672 129 2792 173
rect 2896 129 3016 173
rect 3064 81 3184 173
rect 132 25 252 69
rect 356 25 476 69
rect 624 41 3184 81
rect 3328 25 3448 69
rect 3552 25 3672 69
<< polycontact >>
rect 417 366 463 412
rect 685 477 731 523
rect 1021 384 1067 430
rect 1225 494 1271 540
rect 1889 384 1935 430
rect 2724 366 2770 412
rect 2942 441 2988 487
rect 3341 366 3387 508
<< metal1 >>
rect 0 920 3808 1098
rect 0 918 121 920
rect 167 918 529 920
rect 121 769 167 780
rect 575 918 3637 920
rect 1557 838 1603 918
rect 1557 781 1603 792
rect 2005 838 2051 918
rect 529 769 575 780
rect 254 726 371 766
rect 1761 737 1807 748
rect 254 586 325 726
rect 1109 726 1155 737
rect 254 320 371 586
rect 593 588 1109 634
rect 593 423 639 588
rect 1342 586 1353 632
rect 1399 597 1761 632
rect 2353 838 2399 918
rect 2005 687 2051 698
rect 2149 737 2195 748
rect 1399 586 1807 597
rect 3193 838 3239 918
rect 3193 781 3239 792
rect 3683 918 3808 920
rect 3637 769 3683 780
rect 2353 687 2399 698
rect 2577 737 2623 748
rect 2195 597 2577 632
rect 3433 726 3479 737
rect 2149 586 2623 597
rect 2821 632 3387 643
rect 2867 597 3387 632
rect 1109 575 1155 586
rect 685 523 921 542
rect 2821 540 2867 586
rect 731 477 921 523
rect 1214 494 1225 540
rect 1271 494 2867 540
rect 685 466 921 477
rect 2942 487 3222 542
rect 2988 441 3222 487
rect 2942 430 3222 441
rect 3341 508 3387 597
rect 417 412 639 423
rect 463 366 639 412
rect 1010 384 1021 430
rect 1067 384 1889 430
rect 1935 412 2770 430
rect 1935 384 2724 412
rect 417 355 639 366
rect 57 222 103 233
rect 0 82 57 90
rect 254 180 281 320
rect 327 180 371 320
rect 593 320 639 355
rect 2718 366 2724 384
rect 2718 354 2770 366
rect 1333 320 1827 335
rect 593 274 1109 320
rect 1155 274 1166 320
rect 1379 289 1781 320
rect 1333 263 1379 274
rect 1781 263 1827 274
rect 2149 320 2643 335
rect 3341 331 3387 366
rect 2195 289 2597 320
rect 2149 263 2195 274
rect 2810 320 3387 331
rect 2810 274 2821 320
rect 2867 285 3387 320
rect 3433 542 3479 586
rect 3433 320 3554 542
rect 2867 274 2878 285
rect 2597 263 2643 274
rect 254 169 371 180
rect 505 222 551 233
rect 103 82 505 90
rect 1557 232 1603 243
rect 1557 90 1603 186
rect 2005 232 2051 243
rect 2005 90 2051 186
rect 2373 232 2419 243
rect 2373 90 2419 186
rect 3253 228 3299 239
rect 3253 90 3299 182
rect 3433 180 3477 320
rect 3523 180 3554 320
rect 3433 169 3554 180
rect 3701 222 3747 233
rect 551 82 3701 90
rect 3747 82 3808 90
rect 0 -90 3808 82
<< labels >>
flabel metal1 s 685 466 921 542 0 FreeSans 200 0 0 0 A
port 1 nsew default input
flabel metal1 s 2942 430 3222 542 0 FreeSans 200 0 0 0 B
port 2 nsew default input
flabel metal1 s 1010 384 2770 430 0 FreeSans 200 0 0 0 CI
port 3 nsew default input
flabel metal1 s 3433 542 3479 737 0 FreeSans 200 0 0 0 CO
port 4 nsew default output
flabel metal1 s 254 169 371 766 0 FreeSans 200 0 0 0 S
port 5 nsew default output
flabel metal1 s 0 918 3808 1098 0 FreeSans 200 0 0 0 VDD
port 6 nsew power bidirectional abutment
flabel metal1 s 2373 239 2419 243 0 FreeSans 200 0 0 0 VSS
port 9 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 2718 354 2770 384 1 CI
port 3 nsew default input
rlabel metal1 s 3433 169 3554 542 1 CO
port 4 nsew default output
rlabel metal1 s 3637 781 3683 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3193 781 3239 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2353 781 2399 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2005 781 2051 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 1557 781 1603 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 529 781 575 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 121 781 167 918 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 3637 769 3683 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2353 769 2399 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2005 769 2051 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 529 769 575 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 121 769 167 781 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2353 687 2399 769 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2005 687 2051 769 1 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 2005 239 2051 243 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1557 239 1603 243 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3253 233 3299 239 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2373 233 2419 239 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2005 233 2051 239 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1557 233 1603 239 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3701 90 3747 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 3253 90 3299 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2373 90 2419 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 2005 90 2051 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 1557 90 1603 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 505 90 551 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 57 90 103 233 1 VSS
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3808 90 1 VSS
port 7 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3808 1008
string GDS_END 1073118
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1065358
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
