magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -169 355 170 393
rect -169 299 -134 355
rect -78 299 78 355
rect 134 299 170 355
rect -169 137 170 299
rect -169 81 -134 137
rect -78 81 78 137
rect 134 81 170 137
rect -169 -81 170 81
rect -169 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 170 -81
rect -169 -299 170 -137
rect -169 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 170 -299
rect -169 -393 170 -355
<< via2 >>
rect -134 299 -78 355
rect 78 299 134 355
rect -134 81 -78 137
rect 78 81 134 137
rect -134 -137 -78 -81
rect 78 -137 134 -81
rect -134 -355 -78 -299
rect 78 -355 134 -299
<< metal3 >>
rect -170 355 170 393
rect -170 299 -134 355
rect -78 299 78 355
rect 134 299 170 355
rect -170 137 170 299
rect -170 81 -134 137
rect -78 81 78 137
rect 134 81 170 137
rect -170 -81 170 81
rect -170 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 170 -81
rect -170 -299 170 -137
rect -170 -355 -134 -299
rect -78 -355 78 -299
rect 134 -355 170 -299
rect -170 -393 170 -355
<< properties >>
string GDS_END 674112
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 673468
<< end >>
