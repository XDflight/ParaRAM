magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -220 224 1960 228
rect -221 -717 1960 224
<< nsubdiff >>
rect -78 23 1817 80
rect -78 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1817 23
rect -78 -140 1817 -23
rect -78 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1242 -140
rect 1288 -186 1400 -140
rect 1446 -186 1558 -140
rect 1604 -186 1716 -140
rect 1762 -186 1817 -140
rect -78 -304 1817 -186
rect -78 -350 -23 -304
rect 23 -350 135 -304
rect 181 -350 293 -304
rect 339 -350 451 -304
rect 497 -350 610 -304
rect 656 -350 768 -304
rect 814 -350 926 -304
rect 972 -350 1084 -304
rect 1130 -350 1242 -304
rect 1288 -350 1400 -304
rect 1446 -350 1558 -304
rect 1604 -350 1716 -304
rect 1762 -350 1817 -304
rect -78 -467 1817 -350
rect -78 -513 -23 -467
rect 23 -513 135 -467
rect 181 -513 293 -467
rect 339 -513 451 -467
rect 497 -513 610 -467
rect 656 -513 768 -467
rect 814 -513 926 -467
rect 972 -513 1084 -467
rect 1130 -513 1242 -467
rect 1288 -513 1400 -467
rect 1446 -513 1558 -467
rect 1604 -513 1716 -467
rect 1762 -513 1817 -467
rect -78 -570 1817 -513
<< nsubdiffcont >>
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect 1242 -23 1288 23
rect 1400 -23 1446 23
rect 1558 -23 1604 23
rect 1716 -23 1762 23
rect -23 -186 23 -140
rect 135 -186 181 -140
rect 293 -186 339 -140
rect 451 -186 497 -140
rect 610 -186 656 -140
rect 768 -186 814 -140
rect 926 -186 972 -140
rect 1084 -186 1130 -140
rect 1242 -186 1288 -140
rect 1400 -186 1446 -140
rect 1558 -186 1604 -140
rect 1716 -186 1762 -140
rect -23 -350 23 -304
rect 135 -350 181 -304
rect 293 -350 339 -304
rect 451 -350 497 -304
rect 610 -350 656 -304
rect 768 -350 814 -304
rect 926 -350 972 -304
rect 1084 -350 1130 -304
rect 1242 -350 1288 -304
rect 1400 -350 1446 -304
rect 1558 -350 1604 -304
rect 1716 -350 1762 -304
rect -23 -513 23 -467
rect 135 -513 181 -467
rect 293 -513 339 -467
rect 451 -513 497 -467
rect 610 -513 656 -467
rect 768 -513 814 -467
rect 926 -513 972 -467
rect 1084 -513 1130 -467
rect 1242 -513 1288 -467
rect 1400 -513 1446 -467
rect 1558 -513 1604 -467
rect 1716 -513 1762 -467
<< metal1 >>
rect -58 23 1797 60
rect -58 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1797 23
rect -58 -140 1797 -23
rect -58 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1242 -140
rect 1288 -186 1400 -140
rect 1446 -186 1558 -140
rect 1604 -186 1716 -140
rect 1762 -186 1797 -140
rect -58 -304 1797 -186
rect -58 -350 -23 -304
rect 23 -350 135 -304
rect 181 -350 293 -304
rect 339 -350 451 -304
rect 497 -350 610 -304
rect 656 -350 768 -304
rect 814 -350 926 -304
rect 972 -350 1084 -304
rect 1130 -350 1242 -304
rect 1288 -350 1400 -304
rect 1446 -350 1558 -304
rect 1604 -350 1716 -304
rect 1762 -350 1797 -304
rect -58 -467 1797 -350
rect -58 -513 -23 -467
rect 23 -513 135 -467
rect 181 -513 293 -467
rect 339 -513 451 -467
rect 497 -513 610 -467
rect 656 -513 768 -467
rect 814 -513 926 -467
rect 972 -513 1084 -467
rect 1130 -513 1242 -467
rect 1288 -513 1400 -467
rect 1446 -513 1558 -467
rect 1604 -513 1716 -467
rect 1762 -513 1797 -467
rect -58 -550 1797 -513
<< properties >>
string GDS_END 1219350
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1216002
<< end >>
