magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -83 1281 857 2575
rect 1197 1281 2795 2575
<< mvnmos >>
rect 316 354 456 654
rect 1561 354 1701 654
rect 1805 354 1945 654
rect 2049 354 2189 654
rect 2293 354 2433 654
<< mvpmos >>
rect 316 1486 456 2086
rect 1561 1622 1701 2222
rect 1805 1622 1945 2222
rect 2049 1622 2189 2222
rect 2293 1622 2433 2222
<< mvndiff >>
rect 228 641 316 654
rect 228 595 241 641
rect 287 595 316 641
rect 228 527 316 595
rect 228 481 241 527
rect 287 481 316 527
rect 228 413 316 481
rect 228 367 241 413
rect 287 367 316 413
rect 228 354 316 367
rect 456 641 544 654
rect 456 595 485 641
rect 531 595 544 641
rect 456 527 544 595
rect 456 481 485 527
rect 531 481 544 527
rect 456 413 544 481
rect 456 367 485 413
rect 531 367 544 413
rect 456 354 544 367
rect 1473 641 1561 654
rect 1473 595 1486 641
rect 1532 595 1561 641
rect 1473 527 1561 595
rect 1473 481 1486 527
rect 1532 481 1561 527
rect 1473 413 1561 481
rect 1473 367 1486 413
rect 1532 367 1561 413
rect 1473 354 1561 367
rect 1701 641 1805 654
rect 1701 595 1730 641
rect 1776 595 1805 641
rect 1701 527 1805 595
rect 1701 481 1730 527
rect 1776 481 1805 527
rect 1701 413 1805 481
rect 1701 367 1730 413
rect 1776 367 1805 413
rect 1701 354 1805 367
rect 1945 641 2049 654
rect 1945 595 1974 641
rect 2020 595 2049 641
rect 1945 527 2049 595
rect 1945 481 1974 527
rect 2020 481 2049 527
rect 1945 413 2049 481
rect 1945 367 1974 413
rect 2020 367 2049 413
rect 1945 354 2049 367
rect 2189 641 2293 654
rect 2189 595 2218 641
rect 2264 595 2293 641
rect 2189 527 2293 595
rect 2189 481 2218 527
rect 2264 481 2293 527
rect 2189 413 2293 481
rect 2189 367 2218 413
rect 2264 367 2293 413
rect 2189 354 2293 367
rect 2433 641 2521 654
rect 2433 595 2462 641
rect 2508 595 2521 641
rect 2433 527 2521 595
rect 2433 481 2462 527
rect 2508 481 2521 527
rect 2433 413 2521 481
rect 2433 367 2462 413
rect 2508 367 2521 413
rect 2433 354 2521 367
<< mvpdiff >>
rect 228 2073 316 2086
rect 228 2027 241 2073
rect 287 2027 316 2073
rect 228 1968 316 2027
rect 228 1922 241 1968
rect 287 1922 316 1968
rect 228 1863 316 1922
rect 228 1817 241 1863
rect 287 1817 316 1863
rect 228 1757 316 1817
rect 228 1711 241 1757
rect 287 1711 316 1757
rect 228 1651 316 1711
rect 228 1605 241 1651
rect 287 1605 316 1651
rect 228 1545 316 1605
rect 228 1499 241 1545
rect 287 1499 316 1545
rect 228 1486 316 1499
rect 456 2073 544 2086
rect 456 2027 485 2073
rect 531 2027 544 2073
rect 456 1968 544 2027
rect 456 1922 485 1968
rect 531 1922 544 1968
rect 456 1863 544 1922
rect 456 1817 485 1863
rect 531 1817 544 1863
rect 456 1757 544 1817
rect 456 1711 485 1757
rect 531 1711 544 1757
rect 456 1651 544 1711
rect 456 1605 485 1651
rect 531 1605 544 1651
rect 456 1545 544 1605
rect 456 1499 485 1545
rect 531 1499 544 1545
rect 456 1486 544 1499
rect 1473 2209 1561 2222
rect 1473 2163 1486 2209
rect 1532 2163 1561 2209
rect 1473 2104 1561 2163
rect 1473 2058 1486 2104
rect 1532 2058 1561 2104
rect 1473 1999 1561 2058
rect 1473 1953 1486 1999
rect 1532 1953 1561 1999
rect 1473 1893 1561 1953
rect 1473 1847 1486 1893
rect 1532 1847 1561 1893
rect 1473 1787 1561 1847
rect 1473 1741 1486 1787
rect 1532 1741 1561 1787
rect 1473 1681 1561 1741
rect 1473 1635 1486 1681
rect 1532 1635 1561 1681
rect 1473 1622 1561 1635
rect 1701 2209 1805 2222
rect 1701 2163 1730 2209
rect 1776 2163 1805 2209
rect 1701 2104 1805 2163
rect 1701 2058 1730 2104
rect 1776 2058 1805 2104
rect 1701 1999 1805 2058
rect 1701 1953 1730 1999
rect 1776 1953 1805 1999
rect 1701 1893 1805 1953
rect 1701 1847 1730 1893
rect 1776 1847 1805 1893
rect 1701 1787 1805 1847
rect 1701 1741 1730 1787
rect 1776 1741 1805 1787
rect 1701 1681 1805 1741
rect 1701 1635 1730 1681
rect 1776 1635 1805 1681
rect 1701 1622 1805 1635
rect 1945 2209 2049 2222
rect 1945 2163 1974 2209
rect 2020 2163 2049 2209
rect 1945 2104 2049 2163
rect 1945 2058 1974 2104
rect 2020 2058 2049 2104
rect 1945 1999 2049 2058
rect 1945 1953 1974 1999
rect 2020 1953 2049 1999
rect 1945 1893 2049 1953
rect 1945 1847 1974 1893
rect 2020 1847 2049 1893
rect 1945 1787 2049 1847
rect 1945 1741 1974 1787
rect 2020 1741 2049 1787
rect 1945 1681 2049 1741
rect 1945 1635 1974 1681
rect 2020 1635 2049 1681
rect 1945 1622 2049 1635
rect 2189 2209 2293 2222
rect 2189 2163 2218 2209
rect 2264 2163 2293 2209
rect 2189 2104 2293 2163
rect 2189 2058 2218 2104
rect 2264 2058 2293 2104
rect 2189 1999 2293 2058
rect 2189 1953 2218 1999
rect 2264 1953 2293 1999
rect 2189 1893 2293 1953
rect 2189 1847 2218 1893
rect 2264 1847 2293 1893
rect 2189 1787 2293 1847
rect 2189 1741 2218 1787
rect 2264 1741 2293 1787
rect 2189 1681 2293 1741
rect 2189 1635 2218 1681
rect 2264 1635 2293 1681
rect 2189 1622 2293 1635
rect 2433 2209 2521 2222
rect 2433 2163 2462 2209
rect 2508 2163 2521 2209
rect 2433 2104 2521 2163
rect 2433 2058 2462 2104
rect 2508 2058 2521 2104
rect 2433 1999 2521 2058
rect 2433 1953 2462 1999
rect 2508 1953 2521 1999
rect 2433 1893 2521 1953
rect 2433 1847 2462 1893
rect 2508 1847 2521 1893
rect 2433 1787 2521 1847
rect 2433 1741 2462 1787
rect 2508 1741 2521 1787
rect 2433 1681 2521 1741
rect 2433 1635 2462 1681
rect 2508 1635 2521 1681
rect 2433 1622 2521 1635
<< mvndiffc >>
rect 241 595 287 641
rect 241 481 287 527
rect 241 367 287 413
rect 485 595 531 641
rect 485 481 531 527
rect 485 367 531 413
rect 1486 595 1532 641
rect 1486 481 1532 527
rect 1486 367 1532 413
rect 1730 595 1776 641
rect 1730 481 1776 527
rect 1730 367 1776 413
rect 1974 595 2020 641
rect 1974 481 2020 527
rect 1974 367 2020 413
rect 2218 595 2264 641
rect 2218 481 2264 527
rect 2218 367 2264 413
rect 2462 595 2508 641
rect 2462 481 2508 527
rect 2462 367 2508 413
<< mvpdiffc >>
rect 241 2027 287 2073
rect 241 1922 287 1968
rect 241 1817 287 1863
rect 241 1711 287 1757
rect 241 1605 287 1651
rect 241 1499 287 1545
rect 485 2027 531 2073
rect 485 1922 531 1968
rect 485 1817 531 1863
rect 485 1711 531 1757
rect 485 1605 531 1651
rect 485 1499 531 1545
rect 1486 2163 1532 2209
rect 1486 2058 1532 2104
rect 1486 1953 1532 1999
rect 1486 1847 1532 1893
rect 1486 1741 1532 1787
rect 1486 1635 1532 1681
rect 1730 2163 1776 2209
rect 1730 2058 1776 2104
rect 1730 1953 1776 1999
rect 1730 1847 1776 1893
rect 1730 1741 1776 1787
rect 1730 1635 1776 1681
rect 1974 2163 2020 2209
rect 1974 2058 2020 2104
rect 1974 1953 2020 1999
rect 1974 1847 2020 1893
rect 1974 1741 2020 1787
rect 1974 1635 2020 1681
rect 2218 2163 2264 2209
rect 2218 2058 2264 2104
rect 2218 1953 2264 1999
rect 2218 1847 2264 1893
rect 2218 1741 2264 1787
rect 2218 1635 2264 1681
rect 2462 2163 2508 2209
rect 2462 2058 2508 2104
rect 2462 1953 2508 1999
rect 2462 1847 2508 1893
rect 2462 1741 2508 1787
rect 2462 1635 2508 1681
<< psubdiff >>
rect 0 1008 90 1030
rect 0 22 22 1008
rect 68 90 90 1008
rect 684 914 774 936
rect 684 90 706 914
rect 68 68 706 90
rect 68 22 176 68
rect 598 22 706 68
rect 752 22 774 914
rect 0 0 774 22
rect 1280 914 1370 936
rect 1280 22 1302 914
rect 1348 90 1370 914
rect 2622 1008 2712 1030
rect 2622 90 2644 1008
rect 1348 68 2644 90
rect 1348 22 1456 68
rect 2536 22 2644 68
rect 2690 22 2712 1008
rect 1280 0 2712 22
<< nsubdiff >>
rect 0 2470 774 2492
rect 0 1484 22 2470
rect 68 2424 176 2470
rect 598 2424 706 2470
rect 68 2402 706 2424
rect 68 1484 90 2402
rect 0 1462 90 1484
rect 684 1484 706 2402
rect 752 1484 774 2470
rect 684 1462 774 1484
rect 1280 2470 2712 2492
rect 1280 1484 1302 2470
rect 1348 2424 1456 2470
rect 2536 2424 2644 2470
rect 1348 2402 2644 2424
rect 1348 1484 1370 2402
rect 1280 1462 1370 1484
rect 2622 1484 2644 2402
rect 2690 1484 2712 2470
rect 2622 1462 2712 1484
<< psubdiffcont >>
rect 22 22 68 1008
rect 176 22 598 68
rect 706 22 752 914
rect 1302 22 1348 914
rect 1456 22 2536 68
rect 2644 22 2690 1008
<< nsubdiffcont >>
rect 22 1484 68 2470
rect 176 2424 598 2470
rect 706 1484 752 2470
rect 1302 1484 1348 2470
rect 1456 2424 2536 2470
rect 2644 1484 2690 2470
<< polysilicon >>
rect 316 2086 456 2130
rect 316 1167 456 1486
rect 1561 2222 1701 2266
rect 1805 2222 1945 2266
rect 2049 2222 2189 2266
rect 2293 2222 2433 2266
rect 316 1027 353 1167
rect 399 1027 456 1167
rect 316 654 456 1027
rect 1561 1202 1701 1622
rect 1805 1202 1945 1622
rect 1561 1167 1945 1202
rect 1561 1027 1598 1167
rect 1644 1027 1945 1167
rect 1561 991 1945 1027
rect 316 310 456 354
rect 1561 654 1701 991
rect 1805 654 1945 991
rect 2049 1202 2189 1622
rect 2293 1202 2433 1622
rect 2049 1167 2433 1202
rect 2049 1027 2086 1167
rect 2132 1027 2433 1167
rect 2049 991 2433 1027
rect 2049 654 2189 991
rect 2293 654 2433 991
rect 1561 310 1701 354
rect 1805 310 1945 354
rect 2049 310 2189 354
rect 2293 310 2433 354
<< polycontact >>
rect 353 1027 399 1167
rect 1598 1027 1644 1167
rect 2086 1027 2132 1167
<< metal1 >>
rect 11 2470 763 2481
rect 11 1484 22 2470
rect 68 2424 176 2470
rect 598 2424 706 2470
rect 68 2413 706 2424
rect 68 1484 79 2413
rect 226 2073 302 2413
rect 226 2027 241 2073
rect 287 2027 302 2073
rect 226 1968 302 2027
rect 226 1922 241 1968
rect 287 1922 302 1968
rect 226 1863 302 1922
rect 226 1817 241 1863
rect 287 1817 302 1863
rect 226 1757 302 1817
rect 226 1711 241 1757
rect 287 1711 302 1757
rect 226 1651 302 1711
rect 226 1605 241 1651
rect 287 1605 302 1651
rect 226 1545 302 1605
rect 226 1499 241 1545
rect 287 1499 302 1545
rect 226 1486 302 1499
rect 470 2073 546 2086
rect 470 2027 485 2073
rect 531 2027 546 2073
rect 470 1968 546 2027
rect 470 1922 485 1968
rect 531 1922 546 1968
rect 470 1863 546 1922
rect 470 1817 485 1863
rect 531 1817 546 1863
rect 470 1757 546 1817
rect 470 1711 485 1757
rect 531 1711 546 1757
rect 470 1651 546 1711
rect 470 1605 485 1651
rect 531 1605 546 1651
rect 470 1545 546 1605
rect 470 1499 485 1545
rect 531 1499 546 1545
rect 11 1473 79 1484
rect 470 1186 546 1499
rect 695 1484 706 2413
rect 752 1484 763 2470
rect 695 1473 763 1484
rect 1291 2470 2701 2481
rect 1291 1484 1302 2470
rect 1348 2424 1456 2470
rect 2536 2424 2644 2470
rect 1348 2413 2644 2424
rect 1348 1484 1359 2413
rect 1471 2209 1547 2413
rect 1471 2163 1486 2209
rect 1532 2163 1547 2209
rect 1471 2104 1547 2163
rect 1471 2058 1486 2104
rect 1532 2058 1547 2104
rect 1471 1999 1547 2058
rect 1471 1953 1486 1999
rect 1532 1953 1547 1999
rect 1471 1893 1547 1953
rect 1471 1847 1486 1893
rect 1532 1847 1547 1893
rect 1471 1787 1547 1847
rect 1471 1741 1486 1787
rect 1532 1741 1547 1787
rect 1471 1681 1547 1741
rect 1471 1635 1486 1681
rect 1532 1635 1547 1681
rect 1471 1622 1547 1635
rect 1715 2209 1791 2222
rect 1715 2163 1730 2209
rect 1776 2163 1791 2209
rect 1715 2104 1791 2163
rect 1715 2058 1730 2104
rect 1776 2058 1791 2104
rect 1715 1999 1791 2058
rect 1715 1953 1730 1999
rect 1776 1953 1791 1999
rect 1715 1893 1791 1953
rect 1715 1847 1730 1893
rect 1776 1847 1791 1893
rect 1715 1787 1791 1847
rect 1715 1741 1730 1787
rect 1776 1741 1791 1787
rect 1715 1681 1791 1741
rect 1715 1635 1730 1681
rect 1776 1635 1791 1681
rect 1291 1473 1359 1484
rect 1715 1186 1791 1635
rect 1959 2209 2035 2413
rect 1959 2163 1974 2209
rect 2020 2163 2035 2209
rect 1959 2104 2035 2163
rect 1959 2058 1974 2104
rect 2020 2058 2035 2104
rect 1959 1999 2035 2058
rect 1959 1953 1974 1999
rect 2020 1953 2035 1999
rect 1959 1893 2035 1953
rect 1959 1847 1974 1893
rect 2020 1847 2035 1893
rect 1959 1787 2035 1847
rect 1959 1741 1974 1787
rect 2020 1741 2035 1787
rect 1959 1681 2035 1741
rect 1959 1635 1974 1681
rect 2020 1635 2035 1681
rect 1959 1622 2035 1635
rect 2203 2209 2279 2222
rect 2203 2163 2218 2209
rect 2264 2163 2279 2209
rect 2203 2104 2279 2163
rect 2203 2058 2218 2104
rect 2264 2058 2279 2104
rect 2203 1999 2279 2058
rect 2203 1953 2218 1999
rect 2264 1953 2279 1999
rect 2203 1893 2279 1953
rect 2203 1847 2218 1893
rect 2264 1847 2279 1893
rect 2203 1787 2279 1847
rect 2203 1741 2218 1787
rect 2264 1741 2279 1787
rect 2203 1681 2279 1741
rect 2203 1635 2218 1681
rect 2264 1635 2279 1681
rect 342 1167 410 1178
rect 342 1027 353 1167
rect 399 1027 410 1167
rect 11 1008 79 1019
rect 342 1016 410 1027
rect 470 1167 1655 1186
rect 470 1027 1598 1167
rect 1644 1027 1655 1167
rect 11 22 22 1008
rect 68 79 79 1008
rect 470 1008 1655 1027
rect 1715 1167 2143 1186
rect 1715 1027 2086 1167
rect 2132 1027 2143 1167
rect 1715 1008 2143 1027
rect 226 641 302 654
rect 226 595 241 641
rect 287 595 302 641
rect 226 527 302 595
rect 226 481 241 527
rect 287 481 302 527
rect 226 413 302 481
rect 226 367 241 413
rect 287 367 302 413
rect 226 79 302 367
rect 470 641 546 1008
rect 470 595 485 641
rect 531 595 546 641
rect 470 527 546 595
rect 470 481 485 527
rect 531 481 546 527
rect 470 413 546 481
rect 470 367 485 413
rect 531 367 546 413
rect 470 354 546 367
rect 695 914 763 925
rect 695 79 706 914
rect 68 68 706 79
rect 68 22 176 68
rect 598 22 706 68
rect 752 22 763 914
rect 11 11 763 22
rect 1291 914 1359 925
rect 1291 22 1302 914
rect 1348 79 1359 914
rect 1471 641 1547 654
rect 1471 595 1486 641
rect 1532 595 1547 641
rect 1471 527 1547 595
rect 1471 481 1486 527
rect 1532 481 1547 527
rect 1471 413 1547 481
rect 1471 367 1486 413
rect 1532 367 1547 413
rect 1471 79 1547 367
rect 1715 641 1791 1008
rect 1715 595 1730 641
rect 1776 595 1791 641
rect 1715 527 1791 595
rect 1715 481 1730 527
rect 1776 481 1791 527
rect 1715 413 1791 481
rect 1715 367 1730 413
rect 1776 367 1791 413
rect 1715 354 1791 367
rect 1959 641 2035 654
rect 1959 595 1974 641
rect 2020 595 2035 641
rect 1959 527 2035 595
rect 1959 481 1974 527
rect 2020 481 2035 527
rect 1959 413 2035 481
rect 1959 367 1974 413
rect 2020 367 2035 413
rect 1959 79 2035 367
rect 2203 641 2279 1635
rect 2447 2209 2523 2413
rect 2447 2163 2462 2209
rect 2508 2163 2523 2209
rect 2447 2104 2523 2163
rect 2447 2058 2462 2104
rect 2508 2058 2523 2104
rect 2447 1999 2523 2058
rect 2447 1953 2462 1999
rect 2508 1953 2523 1999
rect 2447 1893 2523 1953
rect 2447 1847 2462 1893
rect 2508 1847 2523 1893
rect 2447 1787 2523 1847
rect 2447 1741 2462 1787
rect 2508 1741 2523 1787
rect 2447 1681 2523 1741
rect 2447 1635 2462 1681
rect 2508 1635 2523 1681
rect 2447 1622 2523 1635
rect 2633 1484 2644 2413
rect 2690 1484 2701 2470
rect 2633 1473 2701 1484
rect 2633 1008 2701 1019
rect 2203 595 2218 641
rect 2264 595 2279 641
rect 2203 527 2279 595
rect 2203 481 2218 527
rect 2264 481 2279 527
rect 2203 413 2279 481
rect 2203 367 2218 413
rect 2264 367 2279 413
rect 2203 354 2279 367
rect 2447 641 2523 654
rect 2447 595 2462 641
rect 2508 595 2523 641
rect 2447 527 2523 595
rect 2447 481 2462 527
rect 2508 481 2523 527
rect 2447 413 2523 481
rect 2447 367 2462 413
rect 2508 367 2523 413
rect 2447 79 2523 367
rect 2633 79 2644 1008
rect 1348 68 2644 79
rect 1348 22 1456 68
rect 2536 22 2644 68
rect 2690 22 2701 1008
rect 1291 11 2701 22
use M1_NWELL_CDNS_40661954729394  M1_NWELL_CDNS_40661954729394_0
timestamp 1666464484
transform 1 0 1996 0 1 2447
box 0 0 1 1
use M1_NWELL_CDNS_40661954729411  M1_NWELL_CDNS_40661954729411_0
timestamp 1666464484
transform 1 0 387 0 1 2447
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_0
timestamp 1666464484
transform 1 0 2667 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_1
timestamp 1666464484
transform 1 0 45 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_2
timestamp 1666464484
transform 1 0 729 0 1 1977
box 0 0 1 1
use M1_NWELL_CDNS_40661954729412  M1_NWELL_CDNS_40661954729412_3
timestamp 1666464484
transform 1 0 1325 0 1 1977
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_0
timestamp 1666464484
transform 1 0 2109 0 1 1097
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_1
timestamp 1666464484
transform 1 0 1621 0 1 1097
box 0 0 1 1
use M1_POLY2_CDNS_40661954729415  M1_POLY2_CDNS_40661954729415_2
timestamp 1666464484
transform 1 0 376 0 1 1097
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_0
timestamp 1666464484
transform 1 0 2667 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661954729413  M1_PSUB_CDNS_40661954729413_1
timestamp 1666464484
transform 1 0 45 0 -1 515
box 0 0 1 1
use M1_PSUB_CDNS_40661954729416  M1_PSUB_CDNS_40661954729416_0
timestamp 1666464484
transform 1 0 387 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661954729422  M1_PSUB_CDNS_40661954729422_0
timestamp 1666464484
transform 1 0 1996 0 -1 45
box 0 0 1 1
use M1_PSUB_CDNS_40661954729423  M1_PSUB_CDNS_40661954729423_0
timestamp 1666464484
transform 1 0 1325 0 -1 468
box 0 0 1 1
use M1_PSUB_CDNS_40661954729423  M1_PSUB_CDNS_40661954729423_1
timestamp 1666464484
transform 1 0 729 0 -1 468
box 0 0 1 1
use nmos_6p0_CDNS_406619547298  nmos_6p0_CDNS_406619547298_0
timestamp 1666464484
transform 1 0 316 0 1 354
box 0 0 1 1
use nmos_6p0_CDNS_4066195472926  nmos_6p0_CDNS_4066195472926_0
timestamp 1666464484
transform 1 0 2049 0 1 354
box 0 0 1 1
use nmos_6p0_CDNS_4066195472926  nmos_6p0_CDNS_4066195472926_1
timestamp 1666464484
transform 1 0 1561 0 1 354
box 0 0 1 1
use pmos_6p0_CDNS_4066195472911  pmos_6p0_CDNS_4066195472911_0
timestamp 1666464484
transform 1 0 316 0 1 1486
box 0 0 1 1
use pmos_6p0_CDNS_4066195472925  pmos_6p0_CDNS_4066195472925_0
timestamp 1666464484
transform 1 0 2049 0 1 1622
box 0 0 1 1
use pmos_6p0_CDNS_4066195472925  pmos_6p0_CDNS_4066195472925_1
timestamp 1666464484
transform 1 0 1561 0 1 1622
box 0 0 1 1
<< labels >>
rlabel metal1 s 1987 1098 1987 1098 4 Z
port 1 nsew
rlabel metal1 s 263 45 263 45 4 VSS
port 2 nsew
rlabel metal1 s 2339 45 2339 45 4 DVSS
port 3 nsew
rlabel metal1 s 2348 2452 2348 2452 4 DVDD
port 4 nsew
rlabel metal1 s 376 1098 376 1098 4 A
port 5 nsew
rlabel metal1 s 29 2452 29 2452 4 VDD
port 6 nsew
rlabel metal1 s 2242 1098 2242 1098 4 ZB
port 7 nsew
<< properties >>
string GDS_END 2031376
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2027458
string path 43.825 8.850 43.825 55.550 
<< end >>
