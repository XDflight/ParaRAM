magic
tech gf180mcuB
timestamp 1666464484
<< properties >>
string GDS_END 2194360
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 2192052
<< end >>
