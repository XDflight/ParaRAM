magic
tech gf180mcuA
magscale 1 5
timestamp 1666464484
<< metal2 >>
rect -236 1161 236 1166
rect -236 1133 -231 1161
rect -203 1133 -169 1161
rect -141 1133 -107 1161
rect -79 1133 -45 1161
rect -17 1133 17 1161
rect 45 1133 79 1161
rect 107 1133 141 1161
rect 169 1133 203 1161
rect 231 1133 236 1161
rect -236 1099 236 1133
rect -236 1071 -231 1099
rect -203 1071 -169 1099
rect -141 1071 -107 1099
rect -79 1071 -45 1099
rect -17 1071 17 1099
rect 45 1071 79 1099
rect 107 1071 141 1099
rect 169 1071 203 1099
rect 231 1071 236 1099
rect -236 1037 236 1071
rect -236 1009 -231 1037
rect -203 1009 -169 1037
rect -141 1009 -107 1037
rect -79 1009 -45 1037
rect -17 1009 17 1037
rect 45 1009 79 1037
rect 107 1009 141 1037
rect 169 1009 203 1037
rect 231 1009 236 1037
rect -236 975 236 1009
rect -236 947 -231 975
rect -203 947 -169 975
rect -141 947 -107 975
rect -79 947 -45 975
rect -17 947 17 975
rect 45 947 79 975
rect 107 947 141 975
rect 169 947 203 975
rect 231 947 236 975
rect -236 913 236 947
rect -236 885 -231 913
rect -203 885 -169 913
rect -141 885 -107 913
rect -79 885 -45 913
rect -17 885 17 913
rect 45 885 79 913
rect 107 885 141 913
rect 169 885 203 913
rect 231 885 236 913
rect -236 851 236 885
rect -236 823 -231 851
rect -203 823 -169 851
rect -141 823 -107 851
rect -79 823 -45 851
rect -17 823 17 851
rect 45 823 79 851
rect 107 823 141 851
rect 169 823 203 851
rect 231 823 236 851
rect -236 789 236 823
rect -236 761 -231 789
rect -203 761 -169 789
rect -141 761 -107 789
rect -79 761 -45 789
rect -17 761 17 789
rect 45 761 79 789
rect 107 761 141 789
rect 169 761 203 789
rect 231 761 236 789
rect -236 727 236 761
rect -236 699 -231 727
rect -203 699 -169 727
rect -141 699 -107 727
rect -79 699 -45 727
rect -17 699 17 727
rect 45 699 79 727
rect 107 699 141 727
rect 169 699 203 727
rect 231 699 236 727
rect -236 665 236 699
rect -236 637 -231 665
rect -203 637 -169 665
rect -141 637 -107 665
rect -79 637 -45 665
rect -17 637 17 665
rect 45 637 79 665
rect 107 637 141 665
rect 169 637 203 665
rect 231 637 236 665
rect -236 603 236 637
rect -236 575 -231 603
rect -203 575 -169 603
rect -141 575 -107 603
rect -79 575 -45 603
rect -17 575 17 603
rect 45 575 79 603
rect 107 575 141 603
rect 169 575 203 603
rect 231 575 236 603
rect -236 541 236 575
rect -236 513 -231 541
rect -203 513 -169 541
rect -141 513 -107 541
rect -79 513 -45 541
rect -17 513 17 541
rect 45 513 79 541
rect 107 513 141 541
rect 169 513 203 541
rect 231 513 236 541
rect -236 479 236 513
rect -236 451 -231 479
rect -203 451 -169 479
rect -141 451 -107 479
rect -79 451 -45 479
rect -17 451 17 479
rect 45 451 79 479
rect 107 451 141 479
rect 169 451 203 479
rect 231 451 236 479
rect -236 417 236 451
rect -236 389 -231 417
rect -203 389 -169 417
rect -141 389 -107 417
rect -79 389 -45 417
rect -17 389 17 417
rect 45 389 79 417
rect 107 389 141 417
rect 169 389 203 417
rect 231 389 236 417
rect -236 355 236 389
rect -236 327 -231 355
rect -203 327 -169 355
rect -141 327 -107 355
rect -79 327 -45 355
rect -17 327 17 355
rect 45 327 79 355
rect 107 327 141 355
rect 169 327 203 355
rect 231 327 236 355
rect -236 293 236 327
rect -236 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 236 293
rect -236 231 236 265
rect -236 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 236 231
rect -236 169 236 203
rect -236 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 236 169
rect -236 107 236 141
rect -236 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 236 107
rect -236 45 236 79
rect -236 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 236 45
rect -236 -17 236 17
rect -236 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 236 -17
rect -236 -79 236 -45
rect -236 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 236 -79
rect -236 -141 236 -107
rect -236 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 236 -141
rect -236 -203 236 -169
rect -236 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 236 -203
rect -236 -265 236 -231
rect -236 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 236 -265
rect -236 -327 236 -293
rect -236 -355 -231 -327
rect -203 -355 -169 -327
rect -141 -355 -107 -327
rect -79 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 79 -327
rect 107 -355 141 -327
rect 169 -355 203 -327
rect 231 -355 236 -327
rect -236 -389 236 -355
rect -236 -417 -231 -389
rect -203 -417 -169 -389
rect -141 -417 -107 -389
rect -79 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 79 -389
rect 107 -417 141 -389
rect 169 -417 203 -389
rect 231 -417 236 -389
rect -236 -451 236 -417
rect -236 -479 -231 -451
rect -203 -479 -169 -451
rect -141 -479 -107 -451
rect -79 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 79 -451
rect 107 -479 141 -451
rect 169 -479 203 -451
rect 231 -479 236 -451
rect -236 -513 236 -479
rect -236 -541 -231 -513
rect -203 -541 -169 -513
rect -141 -541 -107 -513
rect -79 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 79 -513
rect 107 -541 141 -513
rect 169 -541 203 -513
rect 231 -541 236 -513
rect -236 -575 236 -541
rect -236 -603 -231 -575
rect -203 -603 -169 -575
rect -141 -603 -107 -575
rect -79 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 79 -575
rect 107 -603 141 -575
rect 169 -603 203 -575
rect 231 -603 236 -575
rect -236 -637 236 -603
rect -236 -665 -231 -637
rect -203 -665 -169 -637
rect -141 -665 -107 -637
rect -79 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 79 -637
rect 107 -665 141 -637
rect 169 -665 203 -637
rect 231 -665 236 -637
rect -236 -699 236 -665
rect -236 -727 -231 -699
rect -203 -727 -169 -699
rect -141 -727 -107 -699
rect -79 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 79 -699
rect 107 -727 141 -699
rect 169 -727 203 -699
rect 231 -727 236 -699
rect -236 -761 236 -727
rect -236 -789 -231 -761
rect -203 -789 -169 -761
rect -141 -789 -107 -761
rect -79 -789 -45 -761
rect -17 -789 17 -761
rect 45 -789 79 -761
rect 107 -789 141 -761
rect 169 -789 203 -761
rect 231 -789 236 -761
rect -236 -823 236 -789
rect -236 -851 -231 -823
rect -203 -851 -169 -823
rect -141 -851 -107 -823
rect -79 -851 -45 -823
rect -17 -851 17 -823
rect 45 -851 79 -823
rect 107 -851 141 -823
rect 169 -851 203 -823
rect 231 -851 236 -823
rect -236 -885 236 -851
rect -236 -913 -231 -885
rect -203 -913 -169 -885
rect -141 -913 -107 -885
rect -79 -913 -45 -885
rect -17 -913 17 -885
rect 45 -913 79 -885
rect 107 -913 141 -885
rect 169 -913 203 -885
rect 231 -913 236 -885
rect -236 -947 236 -913
rect -236 -975 -231 -947
rect -203 -975 -169 -947
rect -141 -975 -107 -947
rect -79 -975 -45 -947
rect -17 -975 17 -947
rect 45 -975 79 -947
rect 107 -975 141 -947
rect 169 -975 203 -947
rect 231 -975 236 -947
rect -236 -1009 236 -975
rect -236 -1037 -231 -1009
rect -203 -1037 -169 -1009
rect -141 -1037 -107 -1009
rect -79 -1037 -45 -1009
rect -17 -1037 17 -1009
rect 45 -1037 79 -1009
rect 107 -1037 141 -1009
rect 169 -1037 203 -1009
rect 231 -1037 236 -1009
rect -236 -1071 236 -1037
rect -236 -1099 -231 -1071
rect -203 -1099 -169 -1071
rect -141 -1099 -107 -1071
rect -79 -1099 -45 -1071
rect -17 -1099 17 -1071
rect 45 -1099 79 -1071
rect 107 -1099 141 -1071
rect 169 -1099 203 -1071
rect 231 -1099 236 -1071
rect -236 -1133 236 -1099
rect -236 -1161 -231 -1133
rect -203 -1161 -169 -1133
rect -141 -1161 -107 -1133
rect -79 -1161 -45 -1133
rect -17 -1161 17 -1133
rect 45 -1161 79 -1133
rect 107 -1161 141 -1133
rect 169 -1161 203 -1133
rect 231 -1161 236 -1133
rect -236 -1166 236 -1161
<< via2 >>
rect -231 1133 -203 1161
rect -169 1133 -141 1161
rect -107 1133 -79 1161
rect -45 1133 -17 1161
rect 17 1133 45 1161
rect 79 1133 107 1161
rect 141 1133 169 1161
rect 203 1133 231 1161
rect -231 1071 -203 1099
rect -169 1071 -141 1099
rect -107 1071 -79 1099
rect -45 1071 -17 1099
rect 17 1071 45 1099
rect 79 1071 107 1099
rect 141 1071 169 1099
rect 203 1071 231 1099
rect -231 1009 -203 1037
rect -169 1009 -141 1037
rect -107 1009 -79 1037
rect -45 1009 -17 1037
rect 17 1009 45 1037
rect 79 1009 107 1037
rect 141 1009 169 1037
rect 203 1009 231 1037
rect -231 947 -203 975
rect -169 947 -141 975
rect -107 947 -79 975
rect -45 947 -17 975
rect 17 947 45 975
rect 79 947 107 975
rect 141 947 169 975
rect 203 947 231 975
rect -231 885 -203 913
rect -169 885 -141 913
rect -107 885 -79 913
rect -45 885 -17 913
rect 17 885 45 913
rect 79 885 107 913
rect 141 885 169 913
rect 203 885 231 913
rect -231 823 -203 851
rect -169 823 -141 851
rect -107 823 -79 851
rect -45 823 -17 851
rect 17 823 45 851
rect 79 823 107 851
rect 141 823 169 851
rect 203 823 231 851
rect -231 761 -203 789
rect -169 761 -141 789
rect -107 761 -79 789
rect -45 761 -17 789
rect 17 761 45 789
rect 79 761 107 789
rect 141 761 169 789
rect 203 761 231 789
rect -231 699 -203 727
rect -169 699 -141 727
rect -107 699 -79 727
rect -45 699 -17 727
rect 17 699 45 727
rect 79 699 107 727
rect 141 699 169 727
rect 203 699 231 727
rect -231 637 -203 665
rect -169 637 -141 665
rect -107 637 -79 665
rect -45 637 -17 665
rect 17 637 45 665
rect 79 637 107 665
rect 141 637 169 665
rect 203 637 231 665
rect -231 575 -203 603
rect -169 575 -141 603
rect -107 575 -79 603
rect -45 575 -17 603
rect 17 575 45 603
rect 79 575 107 603
rect 141 575 169 603
rect 203 575 231 603
rect -231 513 -203 541
rect -169 513 -141 541
rect -107 513 -79 541
rect -45 513 -17 541
rect 17 513 45 541
rect 79 513 107 541
rect 141 513 169 541
rect 203 513 231 541
rect -231 451 -203 479
rect -169 451 -141 479
rect -107 451 -79 479
rect -45 451 -17 479
rect 17 451 45 479
rect 79 451 107 479
rect 141 451 169 479
rect 203 451 231 479
rect -231 389 -203 417
rect -169 389 -141 417
rect -107 389 -79 417
rect -45 389 -17 417
rect 17 389 45 417
rect 79 389 107 417
rect 141 389 169 417
rect 203 389 231 417
rect -231 327 -203 355
rect -169 327 -141 355
rect -107 327 -79 355
rect -45 327 -17 355
rect 17 327 45 355
rect 79 327 107 355
rect 141 327 169 355
rect 203 327 231 355
rect -231 265 -203 293
rect -169 265 -141 293
rect -107 265 -79 293
rect -45 265 -17 293
rect 17 265 45 293
rect 79 265 107 293
rect 141 265 169 293
rect 203 265 231 293
rect -231 203 -203 231
rect -169 203 -141 231
rect -107 203 -79 231
rect -45 203 -17 231
rect 17 203 45 231
rect 79 203 107 231
rect 141 203 169 231
rect 203 203 231 231
rect -231 141 -203 169
rect -169 141 -141 169
rect -107 141 -79 169
rect -45 141 -17 169
rect 17 141 45 169
rect 79 141 107 169
rect 141 141 169 169
rect 203 141 231 169
rect -231 79 -203 107
rect -169 79 -141 107
rect -107 79 -79 107
rect -45 79 -17 107
rect 17 79 45 107
rect 79 79 107 107
rect 141 79 169 107
rect 203 79 231 107
rect -231 17 -203 45
rect -169 17 -141 45
rect -107 17 -79 45
rect -45 17 -17 45
rect 17 17 45 45
rect 79 17 107 45
rect 141 17 169 45
rect 203 17 231 45
rect -231 -45 -203 -17
rect -169 -45 -141 -17
rect -107 -45 -79 -17
rect -45 -45 -17 -17
rect 17 -45 45 -17
rect 79 -45 107 -17
rect 141 -45 169 -17
rect 203 -45 231 -17
rect -231 -107 -203 -79
rect -169 -107 -141 -79
rect -107 -107 -79 -79
rect -45 -107 -17 -79
rect 17 -107 45 -79
rect 79 -107 107 -79
rect 141 -107 169 -79
rect 203 -107 231 -79
rect -231 -169 -203 -141
rect -169 -169 -141 -141
rect -107 -169 -79 -141
rect -45 -169 -17 -141
rect 17 -169 45 -141
rect 79 -169 107 -141
rect 141 -169 169 -141
rect 203 -169 231 -141
rect -231 -231 -203 -203
rect -169 -231 -141 -203
rect -107 -231 -79 -203
rect -45 -231 -17 -203
rect 17 -231 45 -203
rect 79 -231 107 -203
rect 141 -231 169 -203
rect 203 -231 231 -203
rect -231 -293 -203 -265
rect -169 -293 -141 -265
rect -107 -293 -79 -265
rect -45 -293 -17 -265
rect 17 -293 45 -265
rect 79 -293 107 -265
rect 141 -293 169 -265
rect 203 -293 231 -265
rect -231 -355 -203 -327
rect -169 -355 -141 -327
rect -107 -355 -79 -327
rect -45 -355 -17 -327
rect 17 -355 45 -327
rect 79 -355 107 -327
rect 141 -355 169 -327
rect 203 -355 231 -327
rect -231 -417 -203 -389
rect -169 -417 -141 -389
rect -107 -417 -79 -389
rect -45 -417 -17 -389
rect 17 -417 45 -389
rect 79 -417 107 -389
rect 141 -417 169 -389
rect 203 -417 231 -389
rect -231 -479 -203 -451
rect -169 -479 -141 -451
rect -107 -479 -79 -451
rect -45 -479 -17 -451
rect 17 -479 45 -451
rect 79 -479 107 -451
rect 141 -479 169 -451
rect 203 -479 231 -451
rect -231 -541 -203 -513
rect -169 -541 -141 -513
rect -107 -541 -79 -513
rect -45 -541 -17 -513
rect 17 -541 45 -513
rect 79 -541 107 -513
rect 141 -541 169 -513
rect 203 -541 231 -513
rect -231 -603 -203 -575
rect -169 -603 -141 -575
rect -107 -603 -79 -575
rect -45 -603 -17 -575
rect 17 -603 45 -575
rect 79 -603 107 -575
rect 141 -603 169 -575
rect 203 -603 231 -575
rect -231 -665 -203 -637
rect -169 -665 -141 -637
rect -107 -665 -79 -637
rect -45 -665 -17 -637
rect 17 -665 45 -637
rect 79 -665 107 -637
rect 141 -665 169 -637
rect 203 -665 231 -637
rect -231 -727 -203 -699
rect -169 -727 -141 -699
rect -107 -727 -79 -699
rect -45 -727 -17 -699
rect 17 -727 45 -699
rect 79 -727 107 -699
rect 141 -727 169 -699
rect 203 -727 231 -699
rect -231 -789 -203 -761
rect -169 -789 -141 -761
rect -107 -789 -79 -761
rect -45 -789 -17 -761
rect 17 -789 45 -761
rect 79 -789 107 -761
rect 141 -789 169 -761
rect 203 -789 231 -761
rect -231 -851 -203 -823
rect -169 -851 -141 -823
rect -107 -851 -79 -823
rect -45 -851 -17 -823
rect 17 -851 45 -823
rect 79 -851 107 -823
rect 141 -851 169 -823
rect 203 -851 231 -823
rect -231 -913 -203 -885
rect -169 -913 -141 -885
rect -107 -913 -79 -885
rect -45 -913 -17 -885
rect 17 -913 45 -885
rect 79 -913 107 -885
rect 141 -913 169 -885
rect 203 -913 231 -885
rect -231 -975 -203 -947
rect -169 -975 -141 -947
rect -107 -975 -79 -947
rect -45 -975 -17 -947
rect 17 -975 45 -947
rect 79 -975 107 -947
rect 141 -975 169 -947
rect 203 -975 231 -947
rect -231 -1037 -203 -1009
rect -169 -1037 -141 -1009
rect -107 -1037 -79 -1009
rect -45 -1037 -17 -1009
rect 17 -1037 45 -1009
rect 79 -1037 107 -1009
rect 141 -1037 169 -1009
rect 203 -1037 231 -1009
rect -231 -1099 -203 -1071
rect -169 -1099 -141 -1071
rect -107 -1099 -79 -1071
rect -45 -1099 -17 -1071
rect 17 -1099 45 -1071
rect 79 -1099 107 -1071
rect 141 -1099 169 -1071
rect 203 -1099 231 -1071
rect -231 -1161 -203 -1133
rect -169 -1161 -141 -1133
rect -107 -1161 -79 -1133
rect -45 -1161 -17 -1133
rect 17 -1161 45 -1133
rect 79 -1161 107 -1133
rect 141 -1161 169 -1133
rect 203 -1161 231 -1133
<< metal3 >>
rect -236 1161 236 1166
rect -236 1133 -231 1161
rect -203 1133 -169 1161
rect -141 1133 -107 1161
rect -79 1133 -45 1161
rect -17 1133 17 1161
rect 45 1133 79 1161
rect 107 1133 141 1161
rect 169 1133 203 1161
rect 231 1133 236 1161
rect -236 1099 236 1133
rect -236 1071 -231 1099
rect -203 1071 -169 1099
rect -141 1071 -107 1099
rect -79 1071 -45 1099
rect -17 1071 17 1099
rect 45 1071 79 1099
rect 107 1071 141 1099
rect 169 1071 203 1099
rect 231 1071 236 1099
rect -236 1037 236 1071
rect -236 1009 -231 1037
rect -203 1009 -169 1037
rect -141 1009 -107 1037
rect -79 1009 -45 1037
rect -17 1009 17 1037
rect 45 1009 79 1037
rect 107 1009 141 1037
rect 169 1009 203 1037
rect 231 1009 236 1037
rect -236 975 236 1009
rect -236 947 -231 975
rect -203 947 -169 975
rect -141 947 -107 975
rect -79 947 -45 975
rect -17 947 17 975
rect 45 947 79 975
rect 107 947 141 975
rect 169 947 203 975
rect 231 947 236 975
rect -236 913 236 947
rect -236 885 -231 913
rect -203 885 -169 913
rect -141 885 -107 913
rect -79 885 -45 913
rect -17 885 17 913
rect 45 885 79 913
rect 107 885 141 913
rect 169 885 203 913
rect 231 885 236 913
rect -236 851 236 885
rect -236 823 -231 851
rect -203 823 -169 851
rect -141 823 -107 851
rect -79 823 -45 851
rect -17 823 17 851
rect 45 823 79 851
rect 107 823 141 851
rect 169 823 203 851
rect 231 823 236 851
rect -236 789 236 823
rect -236 761 -231 789
rect -203 761 -169 789
rect -141 761 -107 789
rect -79 761 -45 789
rect -17 761 17 789
rect 45 761 79 789
rect 107 761 141 789
rect 169 761 203 789
rect 231 761 236 789
rect -236 727 236 761
rect -236 699 -231 727
rect -203 699 -169 727
rect -141 699 -107 727
rect -79 699 -45 727
rect -17 699 17 727
rect 45 699 79 727
rect 107 699 141 727
rect 169 699 203 727
rect 231 699 236 727
rect -236 665 236 699
rect -236 637 -231 665
rect -203 637 -169 665
rect -141 637 -107 665
rect -79 637 -45 665
rect -17 637 17 665
rect 45 637 79 665
rect 107 637 141 665
rect 169 637 203 665
rect 231 637 236 665
rect -236 603 236 637
rect -236 575 -231 603
rect -203 575 -169 603
rect -141 575 -107 603
rect -79 575 -45 603
rect -17 575 17 603
rect 45 575 79 603
rect 107 575 141 603
rect 169 575 203 603
rect 231 575 236 603
rect -236 541 236 575
rect -236 513 -231 541
rect -203 513 -169 541
rect -141 513 -107 541
rect -79 513 -45 541
rect -17 513 17 541
rect 45 513 79 541
rect 107 513 141 541
rect 169 513 203 541
rect 231 513 236 541
rect -236 479 236 513
rect -236 451 -231 479
rect -203 451 -169 479
rect -141 451 -107 479
rect -79 451 -45 479
rect -17 451 17 479
rect 45 451 79 479
rect 107 451 141 479
rect 169 451 203 479
rect 231 451 236 479
rect -236 417 236 451
rect -236 389 -231 417
rect -203 389 -169 417
rect -141 389 -107 417
rect -79 389 -45 417
rect -17 389 17 417
rect 45 389 79 417
rect 107 389 141 417
rect 169 389 203 417
rect 231 389 236 417
rect -236 355 236 389
rect -236 327 -231 355
rect -203 327 -169 355
rect -141 327 -107 355
rect -79 327 -45 355
rect -17 327 17 355
rect 45 327 79 355
rect 107 327 141 355
rect 169 327 203 355
rect 231 327 236 355
rect -236 293 236 327
rect -236 265 -231 293
rect -203 265 -169 293
rect -141 265 -107 293
rect -79 265 -45 293
rect -17 265 17 293
rect 45 265 79 293
rect 107 265 141 293
rect 169 265 203 293
rect 231 265 236 293
rect -236 231 236 265
rect -236 203 -231 231
rect -203 203 -169 231
rect -141 203 -107 231
rect -79 203 -45 231
rect -17 203 17 231
rect 45 203 79 231
rect 107 203 141 231
rect 169 203 203 231
rect 231 203 236 231
rect -236 169 236 203
rect -236 141 -231 169
rect -203 141 -169 169
rect -141 141 -107 169
rect -79 141 -45 169
rect -17 141 17 169
rect 45 141 79 169
rect 107 141 141 169
rect 169 141 203 169
rect 231 141 236 169
rect -236 107 236 141
rect -236 79 -231 107
rect -203 79 -169 107
rect -141 79 -107 107
rect -79 79 -45 107
rect -17 79 17 107
rect 45 79 79 107
rect 107 79 141 107
rect 169 79 203 107
rect 231 79 236 107
rect -236 45 236 79
rect -236 17 -231 45
rect -203 17 -169 45
rect -141 17 -107 45
rect -79 17 -45 45
rect -17 17 17 45
rect 45 17 79 45
rect 107 17 141 45
rect 169 17 203 45
rect 231 17 236 45
rect -236 -17 236 17
rect -236 -45 -231 -17
rect -203 -45 -169 -17
rect -141 -45 -107 -17
rect -79 -45 -45 -17
rect -17 -45 17 -17
rect 45 -45 79 -17
rect 107 -45 141 -17
rect 169 -45 203 -17
rect 231 -45 236 -17
rect -236 -79 236 -45
rect -236 -107 -231 -79
rect -203 -107 -169 -79
rect -141 -107 -107 -79
rect -79 -107 -45 -79
rect -17 -107 17 -79
rect 45 -107 79 -79
rect 107 -107 141 -79
rect 169 -107 203 -79
rect 231 -107 236 -79
rect -236 -141 236 -107
rect -236 -169 -231 -141
rect -203 -169 -169 -141
rect -141 -169 -107 -141
rect -79 -169 -45 -141
rect -17 -169 17 -141
rect 45 -169 79 -141
rect 107 -169 141 -141
rect 169 -169 203 -141
rect 231 -169 236 -141
rect -236 -203 236 -169
rect -236 -231 -231 -203
rect -203 -231 -169 -203
rect -141 -231 -107 -203
rect -79 -231 -45 -203
rect -17 -231 17 -203
rect 45 -231 79 -203
rect 107 -231 141 -203
rect 169 -231 203 -203
rect 231 -231 236 -203
rect -236 -265 236 -231
rect -236 -293 -231 -265
rect -203 -293 -169 -265
rect -141 -293 -107 -265
rect -79 -293 -45 -265
rect -17 -293 17 -265
rect 45 -293 79 -265
rect 107 -293 141 -265
rect 169 -293 203 -265
rect 231 -293 236 -265
rect -236 -327 236 -293
rect -236 -355 -231 -327
rect -203 -355 -169 -327
rect -141 -355 -107 -327
rect -79 -355 -45 -327
rect -17 -355 17 -327
rect 45 -355 79 -327
rect 107 -355 141 -327
rect 169 -355 203 -327
rect 231 -355 236 -327
rect -236 -389 236 -355
rect -236 -417 -231 -389
rect -203 -417 -169 -389
rect -141 -417 -107 -389
rect -79 -417 -45 -389
rect -17 -417 17 -389
rect 45 -417 79 -389
rect 107 -417 141 -389
rect 169 -417 203 -389
rect 231 -417 236 -389
rect -236 -451 236 -417
rect -236 -479 -231 -451
rect -203 -479 -169 -451
rect -141 -479 -107 -451
rect -79 -479 -45 -451
rect -17 -479 17 -451
rect 45 -479 79 -451
rect 107 -479 141 -451
rect 169 -479 203 -451
rect 231 -479 236 -451
rect -236 -513 236 -479
rect -236 -541 -231 -513
rect -203 -541 -169 -513
rect -141 -541 -107 -513
rect -79 -541 -45 -513
rect -17 -541 17 -513
rect 45 -541 79 -513
rect 107 -541 141 -513
rect 169 -541 203 -513
rect 231 -541 236 -513
rect -236 -575 236 -541
rect -236 -603 -231 -575
rect -203 -603 -169 -575
rect -141 -603 -107 -575
rect -79 -603 -45 -575
rect -17 -603 17 -575
rect 45 -603 79 -575
rect 107 -603 141 -575
rect 169 -603 203 -575
rect 231 -603 236 -575
rect -236 -637 236 -603
rect -236 -665 -231 -637
rect -203 -665 -169 -637
rect -141 -665 -107 -637
rect -79 -665 -45 -637
rect -17 -665 17 -637
rect 45 -665 79 -637
rect 107 -665 141 -637
rect 169 -665 203 -637
rect 231 -665 236 -637
rect -236 -699 236 -665
rect -236 -727 -231 -699
rect -203 -727 -169 -699
rect -141 -727 -107 -699
rect -79 -727 -45 -699
rect -17 -727 17 -699
rect 45 -727 79 -699
rect 107 -727 141 -699
rect 169 -727 203 -699
rect 231 -727 236 -699
rect -236 -761 236 -727
rect -236 -789 -231 -761
rect -203 -789 -169 -761
rect -141 -789 -107 -761
rect -79 -789 -45 -761
rect -17 -789 17 -761
rect 45 -789 79 -761
rect 107 -789 141 -761
rect 169 -789 203 -761
rect 231 -789 236 -761
rect -236 -823 236 -789
rect -236 -851 -231 -823
rect -203 -851 -169 -823
rect -141 -851 -107 -823
rect -79 -851 -45 -823
rect -17 -851 17 -823
rect 45 -851 79 -823
rect 107 -851 141 -823
rect 169 -851 203 -823
rect 231 -851 236 -823
rect -236 -885 236 -851
rect -236 -913 -231 -885
rect -203 -913 -169 -885
rect -141 -913 -107 -885
rect -79 -913 -45 -885
rect -17 -913 17 -885
rect 45 -913 79 -885
rect 107 -913 141 -885
rect 169 -913 203 -885
rect 231 -913 236 -885
rect -236 -947 236 -913
rect -236 -975 -231 -947
rect -203 -975 -169 -947
rect -141 -975 -107 -947
rect -79 -975 -45 -947
rect -17 -975 17 -947
rect 45 -975 79 -947
rect 107 -975 141 -947
rect 169 -975 203 -947
rect 231 -975 236 -947
rect -236 -1009 236 -975
rect -236 -1037 -231 -1009
rect -203 -1037 -169 -1009
rect -141 -1037 -107 -1009
rect -79 -1037 -45 -1009
rect -17 -1037 17 -1009
rect 45 -1037 79 -1009
rect 107 -1037 141 -1009
rect 169 -1037 203 -1009
rect 231 -1037 236 -1009
rect -236 -1071 236 -1037
rect -236 -1099 -231 -1071
rect -203 -1099 -169 -1071
rect -141 -1099 -107 -1071
rect -79 -1099 -45 -1071
rect -17 -1099 17 -1071
rect 45 -1099 79 -1071
rect 107 -1099 141 -1071
rect 169 -1099 203 -1071
rect 231 -1099 236 -1071
rect -236 -1133 236 -1099
rect -236 -1161 -231 -1133
rect -203 -1161 -169 -1133
rect -141 -1161 -107 -1133
rect -79 -1161 -45 -1133
rect -17 -1161 17 -1133
rect 45 -1161 79 -1133
rect 107 -1161 141 -1133
rect 169 -1161 203 -1133
rect 231 -1161 236 -1133
rect -236 -1166 236 -1161
<< properties >>
string GDS_END 653980
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 634392
<< end >>
