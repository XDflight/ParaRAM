magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 2662 870
<< pwell >>
rect -86 -86 2662 352
<< mvnmos >>
rect 124 93 244 165
rect 348 93 468 165
rect 608 93 728 165
rect 832 93 952 165
rect 1016 93 1136 165
rect 1387 93 1507 165
rect 1611 93 1731 165
rect 1871 68 1991 232
rect 2095 68 2215 232
rect 2279 68 2399 232
<< mvpmos >>
rect 144 524 244 596
rect 348 524 448 596
rect 618 524 718 637
rect 832 524 932 637
rect 1036 524 1136 637
rect 1424 472 1524 585
rect 1588 472 1688 585
rect 1836 472 1936 716
rect 2040 472 2140 716
rect 2244 472 2344 716
<< mvndiff >>
rect 1791 165 1871 232
rect 36 152 124 165
rect 36 106 49 152
rect 95 106 124 152
rect 36 93 124 106
rect 244 152 348 165
rect 244 106 273 152
rect 319 106 348 152
rect 244 93 348 106
rect 468 152 608 165
rect 468 106 497 152
rect 543 106 608 152
rect 468 93 608 106
rect 728 152 832 165
rect 728 106 757 152
rect 803 106 832 152
rect 728 93 832 106
rect 952 93 1016 165
rect 1136 152 1224 165
rect 1136 106 1165 152
rect 1211 106 1224 152
rect 1136 93 1224 106
rect 1299 152 1387 165
rect 1299 106 1312 152
rect 1358 106 1387 152
rect 1299 93 1387 106
rect 1507 152 1611 165
rect 1507 106 1536 152
rect 1582 106 1611 152
rect 1507 93 1611 106
rect 1731 152 1871 165
rect 1731 106 1796 152
rect 1842 106 1871 152
rect 1731 93 1871 106
rect 1791 68 1871 93
rect 1991 180 2095 232
rect 1991 134 2020 180
rect 2066 134 2095 180
rect 1991 68 2095 134
rect 2215 68 2279 232
rect 2399 127 2487 232
rect 2399 81 2428 127
rect 2474 81 2487 127
rect 2399 68 2487 81
<< mvpdiff >>
rect 1748 703 1836 716
rect 538 596 618 637
rect 56 583 144 596
rect 56 537 69 583
rect 115 537 144 583
rect 56 524 144 537
rect 244 524 348 596
rect 448 583 618 596
rect 448 537 477 583
rect 523 537 618 583
rect 448 524 618 537
rect 718 600 832 637
rect 718 554 757 600
rect 803 554 832 600
rect 718 524 832 554
rect 932 583 1036 637
rect 932 537 961 583
rect 1007 537 1036 583
rect 932 524 1036 537
rect 1136 624 1224 637
rect 1136 578 1165 624
rect 1211 578 1224 624
rect 1748 585 1761 703
rect 1136 524 1224 578
rect 1336 548 1424 585
rect 1336 502 1349 548
rect 1395 502 1424 548
rect 1336 472 1424 502
rect 1524 472 1588 585
rect 1688 563 1761 585
rect 1807 563 1836 703
rect 1688 472 1836 563
rect 1936 678 2040 716
rect 1936 632 1965 678
rect 2011 632 2040 678
rect 1936 472 2040 632
rect 2140 586 2244 716
rect 2140 540 2169 586
rect 2215 540 2244 586
rect 2140 472 2244 540
rect 2344 678 2432 716
rect 2344 632 2373 678
rect 2419 632 2432 678
rect 2344 472 2432 632
<< mvndiffc >>
rect 49 106 95 152
rect 273 106 319 152
rect 497 106 543 152
rect 757 106 803 152
rect 1165 106 1211 152
rect 1312 106 1358 152
rect 1536 106 1582 152
rect 1796 106 1842 152
rect 2020 134 2066 180
rect 2428 81 2474 127
<< mvpdiffc >>
rect 69 537 115 583
rect 477 537 523 583
rect 757 554 803 600
rect 961 537 1007 583
rect 1165 578 1211 624
rect 1349 502 1395 548
rect 1761 563 1807 703
rect 1965 632 2011 678
rect 2169 540 2215 586
rect 2373 632 2419 678
<< polysilicon >>
rect 1836 716 1936 760
rect 2040 716 2140 760
rect 2244 716 2344 760
rect 144 596 244 640
rect 348 596 448 640
rect 618 637 718 681
rect 832 637 932 681
rect 1036 637 1136 681
rect 1424 585 1524 629
rect 1588 585 1688 629
rect 144 470 244 524
rect 144 329 173 470
rect 219 329 244 470
rect 144 209 244 329
rect 124 165 244 209
rect 348 303 448 524
rect 348 257 389 303
rect 435 257 448 303
rect 348 209 448 257
rect 618 399 718 524
rect 618 353 642 399
rect 688 353 718 399
rect 618 209 718 353
rect 832 303 932 524
rect 832 257 858 303
rect 904 257 932 303
rect 832 209 932 257
rect 1036 415 1136 524
rect 1036 369 1059 415
rect 1105 369 1136 415
rect 1036 209 1136 369
rect 1424 276 1524 472
rect 348 165 468 209
rect 608 165 728 209
rect 832 165 952 209
rect 1016 165 1136 209
rect 1387 261 1524 276
rect 1588 352 1688 472
rect 1588 337 1731 352
rect 1588 291 1652 337
rect 1698 291 1731 337
rect 1836 326 1936 472
rect 2040 402 2140 472
rect 2244 415 2344 472
rect 2040 356 2195 402
rect 1836 311 1991 326
rect 1836 292 1891 311
rect 1588 275 1731 291
rect 1387 215 1417 261
rect 1463 225 1524 261
rect 1463 215 1507 225
rect 1387 165 1507 215
rect 1611 165 1731 275
rect 1871 265 1891 292
rect 1937 265 1991 311
rect 1871 232 1991 265
rect 2095 311 2195 356
rect 2244 369 2270 415
rect 2316 369 2344 415
rect 2244 330 2344 369
rect 2095 265 2126 311
rect 2172 288 2195 311
rect 2172 265 2215 288
rect 2095 232 2215 265
rect 2279 276 2344 330
rect 2279 232 2399 276
rect 124 49 244 93
rect 348 49 468 93
rect 608 49 728 93
rect 832 49 952 93
rect 1016 49 1136 93
rect 1387 49 1507 93
rect 1611 49 1731 93
rect 1871 24 1991 68
rect 2095 24 2215 68
rect 2279 24 2399 68
<< polycontact >>
rect 173 329 219 470
rect 389 257 435 303
rect 642 353 688 399
rect 858 257 904 303
rect 1059 369 1105 415
rect 1652 291 1698 337
rect 1417 215 1463 261
rect 1891 265 1937 311
rect 2270 369 2316 415
rect 2126 265 2172 311
<< metal1 >>
rect 0 724 2576 844
rect 69 583 115 596
rect 466 583 534 724
rect 1750 703 1818 724
rect 69 261 115 537
rect 173 491 420 542
rect 466 537 477 583
rect 523 537 534 583
rect 746 632 1211 678
rect 746 600 814 632
rect 746 554 757 600
rect 803 554 814 600
rect 1165 624 1211 632
rect 746 551 814 554
rect 950 537 961 583
rect 1007 537 1018 583
rect 1165 563 1211 578
rect 1257 632 1585 678
rect 950 511 1018 537
rect 1257 511 1303 632
rect 173 470 839 491
rect 219 445 839 470
rect 950 465 1303 511
rect 1349 548 1395 585
rect 783 419 839 445
rect 783 415 1120 419
rect 173 314 219 329
rect 277 353 642 399
rect 688 353 702 399
rect 783 369 1059 415
rect 1105 369 1120 415
rect 783 364 1120 369
rect 277 261 330 353
rect 69 214 330 261
rect 378 303 920 307
rect 378 257 389 303
rect 435 257 858 303
rect 904 257 920 303
rect 1176 261 1222 465
rect 1349 353 1395 502
rect 1539 512 1585 632
rect 1750 563 1761 703
rect 1807 563 1818 703
rect 1928 632 1965 678
rect 2011 632 2373 678
rect 2419 632 2432 678
rect 1750 558 1818 563
rect 2154 540 2169 586
rect 2215 540 2440 586
rect 1539 494 2117 512
rect 1539 466 2317 494
rect 2079 448 2317 466
rect 1641 365 2041 420
rect 1349 307 1586 353
rect 378 253 920 257
rect 262 152 330 214
rect 1039 215 1417 261
rect 1463 215 1478 261
rect 1039 214 1478 215
rect 1525 244 1586 307
rect 1641 337 1709 365
rect 1641 291 1652 337
rect 1698 291 1709 337
rect 1995 312 2041 365
rect 2270 415 2317 448
rect 2316 369 2317 415
rect 2270 352 2317 369
rect 1995 311 2222 312
rect 1879 265 1891 311
rect 1937 265 1949 311
rect 1879 244 1949 265
rect 1995 265 2126 311
rect 2172 265 2222 311
rect 1995 253 2222 265
rect 2376 259 2440 540
rect 1039 152 1085 214
rect 1525 198 1949 244
rect 2312 203 2440 259
rect 2312 200 2366 203
rect 1525 152 1593 198
rect 2009 180 2366 200
rect 38 106 49 152
rect 95 106 106 152
rect 262 106 273 152
rect 319 106 330 152
rect 486 106 497 152
rect 543 106 554 152
rect 740 106 757 152
rect 803 106 1085 152
rect 1154 106 1165 152
rect 1211 106 1312 152
rect 1358 106 1370 152
rect 1525 106 1536 152
rect 1582 106 1593 152
rect 1783 106 1796 152
rect 1842 106 1855 152
rect 2009 134 2020 180
rect 2066 134 2366 180
rect 38 60 106 106
rect 486 60 554 106
rect 1154 60 1370 106
rect 1783 60 1855 106
rect 2417 81 2428 127
rect 2474 81 2485 127
rect 2417 60 2485 81
rect 0 -60 2576 60
<< labels >>
flabel metal1 s 1641 365 2041 420 0 FreeSans 400 0 0 0 A3
port 3 nsew default input
flabel metal1 s 0 724 2576 844 0 FreeSans 400 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 1783 127 1855 152 0 FreeSans 400 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel metal1 s 2154 540 2440 586 0 FreeSans 400 0 0 0 Z
port 4 nsew default output
flabel metal1 s 378 253 920 307 0 FreeSans 400 0 0 0 A1
port 1 nsew default input
flabel metal1 s 173 491 420 542 0 FreeSans 400 0 0 0 A2
port 2 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 173 445 839 491 1 A2
port 2 nsew default input
rlabel metal1 s 783 419 839 445 1 A2
port 2 nsew default input
rlabel metal1 s 173 419 219 445 1 A2
port 2 nsew default input
rlabel metal1 s 783 364 1120 419 1 A2
port 2 nsew default input
rlabel metal1 s 173 364 219 419 1 A2
port 2 nsew default input
rlabel metal1 s 173 314 219 364 1 A2
port 2 nsew default input
rlabel metal1 s 1995 312 2041 365 1 A3
port 3 nsew default input
rlabel metal1 s 1641 312 1709 365 1 A3
port 3 nsew default input
rlabel metal1 s 1995 291 2222 312 1 A3
port 3 nsew default input
rlabel metal1 s 1641 291 1709 312 1 A3
port 3 nsew default input
rlabel metal1 s 1995 253 2222 291 1 A3
port 3 nsew default input
rlabel metal1 s 2376 259 2440 540 1 Z
port 4 nsew default output
rlabel metal1 s 2312 203 2440 259 1 Z
port 4 nsew default output
rlabel metal1 s 2312 200 2366 203 1 Z
port 4 nsew default output
rlabel metal1 s 2009 134 2366 200 1 Z
port 4 nsew default output
rlabel metal1 s 1750 558 1818 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 558 534 724 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 466 537 534 558 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1154 127 1370 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 127 554 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 127 106 152 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2417 60 2485 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1783 60 1855 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1154 60 1370 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 486 60 554 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 127 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2576 60 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 784
string GDS_END 369730
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 363794
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
