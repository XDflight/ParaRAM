magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 29138 95074 56005 95590
rect 29138 93521 32850 95074
rect 35260 94009 39818 95074
rect 35260 93833 39436 94009
rect 45169 93833 49764 95074
rect 52285 93833 56005 95074
<< pwell >>
rect 1774 94682 24710 94714
rect 1774 35138 24710 35170
<< mvpmos >>
rect 7024 32969 7144 33651
rect 7249 32969 7369 33651
rect 7715 32969 7835 33651
rect 7940 32969 8060 33651
rect 17824 32969 17944 33651
rect 18049 32969 18169 33651
rect 18515 32969 18635 33651
rect 18740 32969 18860 33651
rect 66600 32969 66720 33651
rect 66825 32969 66945 33651
rect 67291 32969 67411 33651
rect 67516 32969 67636 33651
rect 77400 32969 77520 33651
rect 77625 32969 77745 33651
rect 78091 32969 78211 33651
rect 78316 32969 78436 33651
rect 7024 32194 7144 32876
rect 7249 32194 7369 32876
rect 7715 32194 7835 32876
rect 7940 32194 8060 32876
rect 17824 32194 17944 32876
rect 18049 32194 18169 32876
rect 18515 32194 18635 32876
rect 18740 32194 18860 32876
rect 66600 32194 66720 32876
rect 66825 32194 66945 32876
rect 67291 32194 67411 32876
rect 67516 32194 67636 32876
rect 77400 32194 77520 32876
rect 77625 32194 77745 32876
rect 78091 32194 78211 32876
rect 78316 32194 78436 32876
<< mvpsubdiff >>
rect 27743 34155 57329 34639
rect 3139 32969 3273 33651
rect 4378 32969 4512 33651
rect 5616 32969 5750 33651
rect 6855 32969 6918 33651
rect 7475 32969 7609 33651
rect 8166 32969 8229 33651
rect 9334 32969 9468 33651
rect 10572 32969 10706 33651
rect 11811 32969 11945 33651
rect 13939 32969 14073 33651
rect 15178 32969 15312 33651
rect 16416 32969 16550 33651
rect 17655 32969 17718 33651
rect 18275 32969 18409 33651
rect 18966 32969 19029 33651
rect 20134 32969 20268 33651
rect 21372 32969 21506 33651
rect 22611 32969 22745 33651
rect 62715 32969 62849 33651
rect 63954 32969 64088 33651
rect 65192 32969 65326 33651
rect 66431 32969 66494 33651
rect 67051 32969 67185 33651
rect 67742 32969 67805 33651
rect 68910 32969 69044 33651
rect 70148 32969 70282 33651
rect 71387 32969 71521 33651
rect 73515 32969 73649 33651
rect 74754 32969 74888 33651
rect 75992 32969 76126 33651
rect 77231 32969 77294 33651
rect 77851 32969 77985 33651
rect 78542 32969 78605 33651
rect 79710 32969 79844 33651
rect 80948 32969 81082 33651
rect 82187 32969 82321 33651
rect 3139 32194 3273 32876
rect 4378 32194 4512 32876
rect 5616 32194 5750 32876
rect 6855 32194 6918 32876
rect 7475 32194 7609 32876
rect 8166 32194 8229 32876
rect 9334 32194 9468 32876
rect 10572 32194 10706 32876
rect 11811 32194 11945 32876
rect 13939 32194 14073 32876
rect 15178 32194 15312 32876
rect 16416 32194 16550 32876
rect 17655 32194 17718 32876
rect 18275 32194 18409 32876
rect 18966 32194 19029 32876
rect 20134 32194 20268 32876
rect 21372 32194 21506 32876
rect 22611 32194 22745 32876
rect 62715 32194 62849 32876
rect 63954 32194 64088 32876
rect 65192 32194 65326 32876
rect 66431 32194 66494 32876
rect 67051 32194 67185 32876
rect 67742 32194 67805 32876
rect 68910 32194 69044 32876
rect 70148 32194 70282 32876
rect 71387 32194 71521 32876
rect 73515 32194 73649 32876
rect 74754 32194 74888 32876
rect 75992 32194 76126 32876
rect 77231 32194 77294 32876
rect 77851 32194 77985 32876
rect 78542 32194 78605 32876
rect 79710 32194 79844 32876
rect 80948 32194 81082 32876
rect 82187 32194 82321 32876
<< metal1 >>
rect 282 95694 86090 96694
rect 282 1282 1282 95694
rect 25312 94454 26039 95694
rect 27607 94653 29197 95694
rect 34227 94671 35013 95694
rect 40062 94671 40590 95694
rect 43738 94671 44564 95694
rect 27607 94601 27790 94653
rect 27842 94601 28001 94653
rect 28053 94601 28212 94653
rect 28264 94601 28423 94653
rect 28475 94601 28634 94653
rect 28686 94601 28845 94653
rect 28897 94601 29056 94653
rect 29108 94601 29197 94653
rect 27607 92853 29197 94601
rect 50098 94485 50913 95694
rect 55927 94653 57736 95694
rect 55927 94601 56015 94653
rect 56067 94601 56226 94653
rect 56278 94601 56437 94653
rect 56489 94601 56648 94653
rect 56700 94601 56859 94653
rect 56911 94601 57070 94653
rect 57122 94601 57281 94653
rect 57333 94601 57736 94653
rect 27607 92801 27790 92853
rect 27842 92801 28001 92853
rect 28053 92801 28212 92853
rect 28264 92801 28423 92853
rect 28475 92801 28634 92853
rect 28686 92801 28845 92853
rect 28897 92801 29056 92853
rect 29108 92801 29197 92853
rect 27607 91053 29197 92801
rect 27607 91001 27790 91053
rect 27842 91001 28001 91053
rect 28053 91001 28212 91053
rect 28264 91001 28423 91053
rect 28475 91001 28634 91053
rect 28686 91001 28845 91053
rect 28897 91001 29056 91053
rect 29108 91001 29197 91053
rect 27607 89253 29197 91001
rect 27607 89201 27790 89253
rect 27842 89201 28001 89253
rect 28053 89201 28212 89253
rect 28264 89201 28423 89253
rect 28475 89201 28634 89253
rect 28686 89201 28845 89253
rect 28897 89201 29056 89253
rect 29108 89201 29197 89253
rect 27607 87453 29197 89201
rect 27607 87401 27790 87453
rect 27842 87401 28001 87453
rect 28053 87401 28212 87453
rect 28264 87401 28423 87453
rect 28475 87401 28634 87453
rect 28686 87401 28845 87453
rect 28897 87401 29056 87453
rect 29108 87401 29197 87453
rect 27607 85653 29197 87401
rect 27607 85601 27790 85653
rect 27842 85601 28001 85653
rect 28053 85601 28212 85653
rect 28264 85601 28423 85653
rect 28475 85601 28634 85653
rect 28686 85601 28845 85653
rect 28897 85601 29056 85653
rect 29108 85601 29197 85653
rect 27607 83853 29197 85601
rect 27607 83801 27790 83853
rect 27842 83801 28001 83853
rect 28053 83801 28212 83853
rect 28264 83801 28423 83853
rect 28475 83801 28634 83853
rect 28686 83801 28845 83853
rect 28897 83801 29056 83853
rect 29108 83801 29197 83853
rect 27607 82053 29197 83801
rect 27607 82001 27790 82053
rect 27842 82001 28001 82053
rect 28053 82001 28212 82053
rect 28264 82001 28423 82053
rect 28475 82001 28634 82053
rect 28686 82001 28845 82053
rect 28897 82001 29056 82053
rect 29108 82001 29197 82053
rect 27607 80253 29197 82001
rect 27607 80201 27790 80253
rect 27842 80201 28001 80253
rect 28053 80201 28212 80253
rect 28264 80201 28423 80253
rect 28475 80201 28634 80253
rect 28686 80201 28845 80253
rect 28897 80201 29056 80253
rect 29108 80201 29197 80253
rect 27607 78453 29197 80201
rect 27607 78401 27790 78453
rect 27842 78401 28001 78453
rect 28053 78401 28212 78453
rect 28264 78401 28423 78453
rect 28475 78401 28634 78453
rect 28686 78401 28845 78453
rect 28897 78401 29056 78453
rect 29108 78401 29197 78453
rect 27607 76653 29197 78401
rect 27607 76601 27790 76653
rect 27842 76601 28001 76653
rect 28053 76601 28212 76653
rect 28264 76601 28423 76653
rect 28475 76601 28634 76653
rect 28686 76601 28845 76653
rect 28897 76601 29056 76653
rect 29108 76601 29197 76653
rect 27607 74853 29197 76601
rect 27607 74801 27790 74853
rect 27842 74801 28001 74853
rect 28053 74801 28212 74853
rect 28264 74801 28423 74853
rect 28475 74801 28634 74853
rect 28686 74801 28845 74853
rect 28897 74801 29056 74853
rect 29108 74801 29197 74853
rect 27607 73053 29197 74801
rect 27607 73001 27790 73053
rect 27842 73001 28001 73053
rect 28053 73001 28212 73053
rect 28264 73001 28423 73053
rect 28475 73001 28634 73053
rect 28686 73001 28845 73053
rect 28897 73001 29056 73053
rect 29108 73001 29197 73053
rect 27607 71253 29197 73001
rect 27607 71201 27790 71253
rect 27842 71201 28001 71253
rect 28053 71201 28212 71253
rect 28264 71201 28423 71253
rect 28475 71201 28634 71253
rect 28686 71201 28845 71253
rect 28897 71201 29056 71253
rect 29108 71201 29197 71253
rect 27607 69453 29197 71201
rect 27607 69401 27790 69453
rect 27842 69401 28001 69453
rect 28053 69401 28212 69453
rect 28264 69401 28423 69453
rect 28475 69401 28634 69453
rect 28686 69401 28845 69453
rect 28897 69401 29056 69453
rect 29108 69401 29197 69453
rect 27607 67653 29197 69401
rect 27607 67601 27790 67653
rect 27842 67601 28001 67653
rect 28053 67601 28212 67653
rect 28264 67601 28423 67653
rect 28475 67601 28634 67653
rect 28686 67601 28845 67653
rect 28897 67601 29056 67653
rect 29108 67601 29197 67653
rect 27607 65853 29197 67601
rect 27607 65801 27790 65853
rect 27842 65801 28001 65853
rect 28053 65801 28212 65853
rect 28264 65801 28423 65853
rect 28475 65801 28634 65853
rect 28686 65801 28845 65853
rect 28897 65801 29056 65853
rect 29108 65801 29197 65853
rect 27607 64053 29197 65801
rect 27607 64001 27790 64053
rect 27842 64001 28001 64053
rect 28053 64001 28212 64053
rect 28264 64001 28423 64053
rect 28475 64001 28634 64053
rect 28686 64001 28845 64053
rect 28897 64001 29056 64053
rect 29108 64001 29197 64053
rect 27607 62253 29197 64001
rect 27607 62201 27790 62253
rect 27842 62201 28001 62253
rect 28053 62201 28212 62253
rect 28264 62201 28423 62253
rect 28475 62201 28634 62253
rect 28686 62201 28845 62253
rect 28897 62201 29056 62253
rect 29108 62201 29197 62253
rect 27607 60453 29197 62201
rect 27607 60401 27790 60453
rect 27842 60401 28001 60453
rect 28053 60401 28212 60453
rect 28264 60401 28423 60453
rect 28475 60401 28634 60453
rect 28686 60401 28845 60453
rect 28897 60401 29056 60453
rect 29108 60401 29197 60453
rect 27607 58653 29197 60401
rect 27607 58601 27790 58653
rect 27842 58601 28001 58653
rect 28053 58601 28212 58653
rect 28264 58601 28423 58653
rect 28475 58601 28634 58653
rect 28686 58601 28845 58653
rect 28897 58601 29056 58653
rect 29108 58601 29197 58653
rect 27607 56853 29197 58601
rect 27607 56801 27790 56853
rect 27842 56801 28001 56853
rect 28053 56801 28212 56853
rect 28264 56801 28423 56853
rect 28475 56801 28634 56853
rect 28686 56801 28845 56853
rect 28897 56801 29056 56853
rect 29108 56801 29197 56853
rect 27607 55053 29197 56801
rect 27607 55001 27790 55053
rect 27842 55001 28001 55053
rect 28053 55001 28212 55053
rect 28264 55001 28423 55053
rect 28475 55001 28634 55053
rect 28686 55001 28845 55053
rect 28897 55001 29056 55053
rect 29108 55001 29197 55053
rect 27607 53253 29197 55001
rect 27607 53201 27790 53253
rect 27842 53201 28001 53253
rect 28053 53201 28212 53253
rect 28264 53201 28423 53253
rect 28475 53201 28634 53253
rect 28686 53201 28845 53253
rect 28897 53201 29056 53253
rect 29108 53201 29197 53253
rect 27607 51453 29197 53201
rect 27607 51401 27790 51453
rect 27842 51401 28001 51453
rect 28053 51401 28212 51453
rect 28264 51401 28423 51453
rect 28475 51401 28634 51453
rect 28686 51401 28845 51453
rect 28897 51401 29056 51453
rect 29108 51401 29197 51453
rect 27607 49653 29197 51401
rect 27607 49601 27790 49653
rect 27842 49601 28001 49653
rect 28053 49601 28212 49653
rect 28264 49601 28423 49653
rect 28475 49601 28634 49653
rect 28686 49601 28845 49653
rect 28897 49601 29056 49653
rect 29108 49601 29197 49653
rect 27607 47853 29197 49601
rect 27607 47801 27790 47853
rect 27842 47801 28001 47853
rect 28053 47801 28212 47853
rect 28264 47801 28423 47853
rect 28475 47801 28634 47853
rect 28686 47801 28845 47853
rect 28897 47801 29056 47853
rect 29108 47801 29197 47853
rect 27607 46053 29197 47801
rect 27607 46001 27790 46053
rect 27842 46001 28001 46053
rect 28053 46001 28212 46053
rect 28264 46001 28423 46053
rect 28475 46001 28634 46053
rect 28686 46001 28845 46053
rect 28897 46001 29056 46053
rect 29108 46001 29197 46053
rect 27607 44253 29197 46001
rect 27607 44201 27790 44253
rect 27842 44201 28001 44253
rect 28053 44201 28212 44253
rect 28264 44201 28423 44253
rect 28475 44201 28634 44253
rect 28686 44201 28845 44253
rect 28897 44201 29056 44253
rect 29108 44201 29197 44253
rect 27607 42453 29197 44201
rect 27607 42401 27790 42453
rect 27842 42401 28001 42453
rect 28053 42401 28212 42453
rect 28264 42401 28423 42453
rect 28475 42401 28634 42453
rect 28686 42401 28845 42453
rect 28897 42401 29056 42453
rect 29108 42401 29197 42453
rect 27607 40653 29197 42401
rect 27607 40601 27790 40653
rect 27842 40601 28001 40653
rect 28053 40601 28212 40653
rect 28264 40601 28423 40653
rect 28475 40601 28634 40653
rect 28686 40601 28845 40653
rect 28897 40601 29056 40653
rect 29108 40601 29197 40653
rect 27607 38853 29197 40601
rect 27607 38801 27790 38853
rect 27842 38801 28001 38853
rect 28053 38801 28212 38853
rect 28264 38801 28423 38853
rect 28475 38801 28634 38853
rect 28686 38801 28845 38853
rect 28897 38801 29056 38853
rect 29108 38801 29197 38853
rect 27607 37053 29197 38801
rect 27607 37001 27790 37053
rect 27842 37001 28001 37053
rect 28053 37001 28212 37053
rect 28264 37001 28423 37053
rect 28475 37001 28634 37053
rect 28686 37001 28845 37053
rect 28897 37001 29056 37053
rect 29108 37001 29197 37053
rect 27607 36421 29197 37001
rect 27387 35985 29197 36421
rect 55927 92853 57736 94601
rect 58791 94454 59518 95694
rect 55927 92801 56015 92853
rect 56067 92801 56226 92853
rect 56278 92801 56437 92853
rect 56489 92801 56648 92853
rect 56700 92801 56859 92853
rect 56911 92801 57070 92853
rect 57122 92801 57281 92853
rect 57333 92801 57736 92853
rect 55927 91053 57736 92801
rect 55927 91001 56015 91053
rect 56067 91001 56226 91053
rect 56278 91001 56437 91053
rect 56489 91001 56648 91053
rect 56700 91001 56859 91053
rect 56911 91001 57070 91053
rect 57122 91001 57281 91053
rect 57333 91001 57736 91053
rect 55927 89253 57736 91001
rect 55927 89201 56015 89253
rect 56067 89201 56226 89253
rect 56278 89201 56437 89253
rect 56489 89201 56648 89253
rect 56700 89201 56859 89253
rect 56911 89201 57070 89253
rect 57122 89201 57281 89253
rect 57333 89201 57736 89253
rect 55927 87453 57736 89201
rect 55927 87401 56015 87453
rect 56067 87401 56226 87453
rect 56278 87401 56437 87453
rect 56489 87401 56648 87453
rect 56700 87401 56859 87453
rect 56911 87401 57070 87453
rect 57122 87401 57281 87453
rect 57333 87401 57736 87453
rect 55927 85653 57736 87401
rect 55927 85601 56015 85653
rect 56067 85601 56226 85653
rect 56278 85601 56437 85653
rect 56489 85601 56648 85653
rect 56700 85601 56859 85653
rect 56911 85601 57070 85653
rect 57122 85601 57281 85653
rect 57333 85601 57736 85653
rect 55927 83853 57736 85601
rect 55927 83801 56015 83853
rect 56067 83801 56226 83853
rect 56278 83801 56437 83853
rect 56489 83801 56648 83853
rect 56700 83801 56859 83853
rect 56911 83801 57070 83853
rect 57122 83801 57281 83853
rect 57333 83801 57736 83853
rect 55927 82053 57736 83801
rect 55927 82001 56015 82053
rect 56067 82001 56226 82053
rect 56278 82001 56437 82053
rect 56489 82001 56648 82053
rect 56700 82001 56859 82053
rect 56911 82001 57070 82053
rect 57122 82001 57281 82053
rect 57333 82001 57736 82053
rect 55927 80253 57736 82001
rect 55927 80201 56015 80253
rect 56067 80201 56226 80253
rect 56278 80201 56437 80253
rect 56489 80201 56648 80253
rect 56700 80201 56859 80253
rect 56911 80201 57070 80253
rect 57122 80201 57281 80253
rect 57333 80201 57736 80253
rect 55927 78453 57736 80201
rect 55927 78401 56015 78453
rect 56067 78401 56226 78453
rect 56278 78401 56437 78453
rect 56489 78401 56648 78453
rect 56700 78401 56859 78453
rect 56911 78401 57070 78453
rect 57122 78401 57281 78453
rect 57333 78401 57736 78453
rect 55927 76653 57736 78401
rect 55927 76601 56015 76653
rect 56067 76601 56226 76653
rect 56278 76601 56437 76653
rect 56489 76601 56648 76653
rect 56700 76601 56859 76653
rect 56911 76601 57070 76653
rect 57122 76601 57281 76653
rect 57333 76601 57736 76653
rect 55927 74853 57736 76601
rect 55927 74801 56015 74853
rect 56067 74801 56226 74853
rect 56278 74801 56437 74853
rect 56489 74801 56648 74853
rect 56700 74801 56859 74853
rect 56911 74801 57070 74853
rect 57122 74801 57281 74853
rect 57333 74801 57736 74853
rect 55927 73053 57736 74801
rect 55927 73001 56015 73053
rect 56067 73001 56226 73053
rect 56278 73001 56437 73053
rect 56489 73001 56648 73053
rect 56700 73001 56859 73053
rect 56911 73001 57070 73053
rect 57122 73001 57281 73053
rect 57333 73001 57736 73053
rect 55927 71253 57736 73001
rect 55927 71201 56015 71253
rect 56067 71201 56226 71253
rect 56278 71201 56437 71253
rect 56489 71201 56648 71253
rect 56700 71201 56859 71253
rect 56911 71201 57070 71253
rect 57122 71201 57281 71253
rect 57333 71201 57736 71253
rect 55927 69453 57736 71201
rect 55927 69401 56015 69453
rect 56067 69401 56226 69453
rect 56278 69401 56437 69453
rect 56489 69401 56648 69453
rect 56700 69401 56859 69453
rect 56911 69401 57070 69453
rect 57122 69401 57281 69453
rect 57333 69401 57736 69453
rect 55927 67653 57736 69401
rect 55927 67601 56015 67653
rect 56067 67601 56226 67653
rect 56278 67601 56437 67653
rect 56489 67601 56648 67653
rect 56700 67601 56859 67653
rect 56911 67601 57070 67653
rect 57122 67601 57281 67653
rect 57333 67601 57736 67653
rect 55927 65853 57736 67601
rect 55927 65801 56015 65853
rect 56067 65801 56226 65853
rect 56278 65801 56437 65853
rect 56489 65801 56648 65853
rect 56700 65801 56859 65853
rect 56911 65801 57070 65853
rect 57122 65801 57281 65853
rect 57333 65801 57736 65853
rect 55927 64053 57736 65801
rect 55927 64001 56015 64053
rect 56067 64001 56226 64053
rect 56278 64001 56437 64053
rect 56489 64001 56648 64053
rect 56700 64001 56859 64053
rect 56911 64001 57070 64053
rect 57122 64001 57281 64053
rect 57333 64001 57736 64053
rect 55927 62253 57736 64001
rect 55927 62201 56015 62253
rect 56067 62201 56226 62253
rect 56278 62201 56437 62253
rect 56489 62201 56648 62253
rect 56700 62201 56859 62253
rect 56911 62201 57070 62253
rect 57122 62201 57281 62253
rect 57333 62201 57736 62253
rect 55927 60453 57736 62201
rect 55927 60401 56015 60453
rect 56067 60401 56226 60453
rect 56278 60401 56437 60453
rect 56489 60401 56648 60453
rect 56700 60401 56859 60453
rect 56911 60401 57070 60453
rect 57122 60401 57281 60453
rect 57333 60401 57736 60453
rect 55927 58653 57736 60401
rect 55927 58601 56015 58653
rect 56067 58601 56226 58653
rect 56278 58601 56437 58653
rect 56489 58601 56648 58653
rect 56700 58601 56859 58653
rect 56911 58601 57070 58653
rect 57122 58601 57281 58653
rect 57333 58601 57736 58653
rect 55927 56853 57736 58601
rect 55927 56801 56015 56853
rect 56067 56801 56226 56853
rect 56278 56801 56437 56853
rect 56489 56801 56648 56853
rect 56700 56801 56859 56853
rect 56911 56801 57070 56853
rect 57122 56801 57281 56853
rect 57333 56801 57736 56853
rect 55927 55053 57736 56801
rect 55927 55001 56015 55053
rect 56067 55001 56226 55053
rect 56278 55001 56437 55053
rect 56489 55001 56648 55053
rect 56700 55001 56859 55053
rect 56911 55001 57070 55053
rect 57122 55001 57281 55053
rect 57333 55001 57736 55053
rect 55927 53253 57736 55001
rect 55927 53201 56015 53253
rect 56067 53201 56226 53253
rect 56278 53201 56437 53253
rect 56489 53201 56648 53253
rect 56700 53201 56859 53253
rect 56911 53201 57070 53253
rect 57122 53201 57281 53253
rect 57333 53201 57736 53253
rect 55927 51453 57736 53201
rect 55927 51401 56015 51453
rect 56067 51401 56226 51453
rect 56278 51401 56437 51453
rect 56489 51401 56648 51453
rect 56700 51401 56859 51453
rect 56911 51401 57070 51453
rect 57122 51401 57281 51453
rect 57333 51401 57736 51453
rect 55927 49653 57736 51401
rect 55927 49601 56015 49653
rect 56067 49601 56226 49653
rect 56278 49601 56437 49653
rect 56489 49601 56648 49653
rect 56700 49601 56859 49653
rect 56911 49601 57070 49653
rect 57122 49601 57281 49653
rect 57333 49601 57736 49653
rect 55927 47853 57736 49601
rect 55927 47801 56015 47853
rect 56067 47801 56226 47853
rect 56278 47801 56437 47853
rect 56489 47801 56648 47853
rect 56700 47801 56859 47853
rect 56911 47801 57070 47853
rect 57122 47801 57281 47853
rect 57333 47801 57736 47853
rect 55927 46053 57736 47801
rect 55927 46001 56015 46053
rect 56067 46001 56226 46053
rect 56278 46001 56437 46053
rect 56489 46001 56648 46053
rect 56700 46001 56859 46053
rect 56911 46001 57070 46053
rect 57122 46001 57281 46053
rect 57333 46001 57736 46053
rect 55927 44253 57736 46001
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44201 56437 44253
rect 56489 44201 56648 44253
rect 56700 44201 56859 44253
rect 56911 44201 57070 44253
rect 57122 44201 57281 44253
rect 57333 44201 57736 44253
rect 55927 42453 57736 44201
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42401 56437 42453
rect 56489 42401 56648 42453
rect 56700 42401 56859 42453
rect 56911 42401 57070 42453
rect 57122 42401 57281 42453
rect 57333 42401 57736 42453
rect 55927 40653 57736 42401
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40601 56437 40653
rect 56489 40601 56648 40653
rect 56700 40601 56859 40653
rect 56911 40601 57070 40653
rect 57122 40601 57281 40653
rect 57333 40601 57736 40653
rect 55927 38853 57736 40601
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38801 56437 38853
rect 56489 38801 56648 38853
rect 56700 38801 56859 38853
rect 56911 38801 57070 38853
rect 57122 38801 57281 38853
rect 57333 38801 57736 38853
rect 55927 37053 57736 38801
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37001 56437 37053
rect 56489 37001 56648 37053
rect 56700 37001 56859 37053
rect 56911 37001 57070 37053
rect 57122 37001 57281 37053
rect 57333 37001 57736 37053
rect 55927 35985 57736 37001
rect 27387 34631 27828 35985
rect 57295 34631 57736 35985
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 85090 35484 86090 95694
rect 84242 35364 86090 35484
rect 60563 35326 60639 35338
rect 27386 34163 57736 34631
rect 26772 1777 27214 33519
rect 27387 1925 27828 34163
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 3584 57736 34163
rect 40611 3282 40791 3294
rect 40611 3230 40623 3282
rect 40779 3230 40791 3282
rect 40611 3218 40791 3230
rect 57295 1925 57737 3584
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1282 57737 1925
rect 57909 1777 58351 33519
rect 83398 32048 83834 32122
rect 62138 1689 62318 1701
rect 62138 1637 62150 1689
rect 62306 1637 62318 1689
rect 62138 1625 62318 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 85090 1282 86090 35364
rect 282 282 86090 1282
<< via1 >>
rect 27790 94601 27842 94653
rect 28001 94601 28053 94653
rect 28212 94601 28264 94653
rect 28423 94601 28475 94653
rect 28634 94601 28686 94653
rect 28845 94601 28897 94653
rect 29056 94601 29108 94653
rect 56015 94601 56067 94653
rect 56226 94601 56278 94653
rect 56437 94601 56489 94653
rect 56648 94601 56700 94653
rect 56859 94601 56911 94653
rect 57070 94601 57122 94653
rect 57281 94601 57333 94653
rect 27790 92801 27842 92853
rect 28001 92801 28053 92853
rect 28212 92801 28264 92853
rect 28423 92801 28475 92853
rect 28634 92801 28686 92853
rect 28845 92801 28897 92853
rect 29056 92801 29108 92853
rect 27790 91001 27842 91053
rect 28001 91001 28053 91053
rect 28212 91001 28264 91053
rect 28423 91001 28475 91053
rect 28634 91001 28686 91053
rect 28845 91001 28897 91053
rect 29056 91001 29108 91053
rect 27790 89201 27842 89253
rect 28001 89201 28053 89253
rect 28212 89201 28264 89253
rect 28423 89201 28475 89253
rect 28634 89201 28686 89253
rect 28845 89201 28897 89253
rect 29056 89201 29108 89253
rect 27790 87401 27842 87453
rect 28001 87401 28053 87453
rect 28212 87401 28264 87453
rect 28423 87401 28475 87453
rect 28634 87401 28686 87453
rect 28845 87401 28897 87453
rect 29056 87401 29108 87453
rect 27790 85601 27842 85653
rect 28001 85601 28053 85653
rect 28212 85601 28264 85653
rect 28423 85601 28475 85653
rect 28634 85601 28686 85653
rect 28845 85601 28897 85653
rect 29056 85601 29108 85653
rect 27790 83801 27842 83853
rect 28001 83801 28053 83853
rect 28212 83801 28264 83853
rect 28423 83801 28475 83853
rect 28634 83801 28686 83853
rect 28845 83801 28897 83853
rect 29056 83801 29108 83853
rect 27790 82001 27842 82053
rect 28001 82001 28053 82053
rect 28212 82001 28264 82053
rect 28423 82001 28475 82053
rect 28634 82001 28686 82053
rect 28845 82001 28897 82053
rect 29056 82001 29108 82053
rect 27790 80201 27842 80253
rect 28001 80201 28053 80253
rect 28212 80201 28264 80253
rect 28423 80201 28475 80253
rect 28634 80201 28686 80253
rect 28845 80201 28897 80253
rect 29056 80201 29108 80253
rect 27790 78401 27842 78453
rect 28001 78401 28053 78453
rect 28212 78401 28264 78453
rect 28423 78401 28475 78453
rect 28634 78401 28686 78453
rect 28845 78401 28897 78453
rect 29056 78401 29108 78453
rect 27790 76601 27842 76653
rect 28001 76601 28053 76653
rect 28212 76601 28264 76653
rect 28423 76601 28475 76653
rect 28634 76601 28686 76653
rect 28845 76601 28897 76653
rect 29056 76601 29108 76653
rect 27790 74801 27842 74853
rect 28001 74801 28053 74853
rect 28212 74801 28264 74853
rect 28423 74801 28475 74853
rect 28634 74801 28686 74853
rect 28845 74801 28897 74853
rect 29056 74801 29108 74853
rect 27790 73001 27842 73053
rect 28001 73001 28053 73053
rect 28212 73001 28264 73053
rect 28423 73001 28475 73053
rect 28634 73001 28686 73053
rect 28845 73001 28897 73053
rect 29056 73001 29108 73053
rect 27790 71201 27842 71253
rect 28001 71201 28053 71253
rect 28212 71201 28264 71253
rect 28423 71201 28475 71253
rect 28634 71201 28686 71253
rect 28845 71201 28897 71253
rect 29056 71201 29108 71253
rect 27790 69401 27842 69453
rect 28001 69401 28053 69453
rect 28212 69401 28264 69453
rect 28423 69401 28475 69453
rect 28634 69401 28686 69453
rect 28845 69401 28897 69453
rect 29056 69401 29108 69453
rect 27790 67601 27842 67653
rect 28001 67601 28053 67653
rect 28212 67601 28264 67653
rect 28423 67601 28475 67653
rect 28634 67601 28686 67653
rect 28845 67601 28897 67653
rect 29056 67601 29108 67653
rect 27790 65801 27842 65853
rect 28001 65801 28053 65853
rect 28212 65801 28264 65853
rect 28423 65801 28475 65853
rect 28634 65801 28686 65853
rect 28845 65801 28897 65853
rect 29056 65801 29108 65853
rect 27790 64001 27842 64053
rect 28001 64001 28053 64053
rect 28212 64001 28264 64053
rect 28423 64001 28475 64053
rect 28634 64001 28686 64053
rect 28845 64001 28897 64053
rect 29056 64001 29108 64053
rect 27790 62201 27842 62253
rect 28001 62201 28053 62253
rect 28212 62201 28264 62253
rect 28423 62201 28475 62253
rect 28634 62201 28686 62253
rect 28845 62201 28897 62253
rect 29056 62201 29108 62253
rect 27790 60401 27842 60453
rect 28001 60401 28053 60453
rect 28212 60401 28264 60453
rect 28423 60401 28475 60453
rect 28634 60401 28686 60453
rect 28845 60401 28897 60453
rect 29056 60401 29108 60453
rect 27790 58601 27842 58653
rect 28001 58601 28053 58653
rect 28212 58601 28264 58653
rect 28423 58601 28475 58653
rect 28634 58601 28686 58653
rect 28845 58601 28897 58653
rect 29056 58601 29108 58653
rect 27790 56801 27842 56853
rect 28001 56801 28053 56853
rect 28212 56801 28264 56853
rect 28423 56801 28475 56853
rect 28634 56801 28686 56853
rect 28845 56801 28897 56853
rect 29056 56801 29108 56853
rect 27790 55001 27842 55053
rect 28001 55001 28053 55053
rect 28212 55001 28264 55053
rect 28423 55001 28475 55053
rect 28634 55001 28686 55053
rect 28845 55001 28897 55053
rect 29056 55001 29108 55053
rect 27790 53201 27842 53253
rect 28001 53201 28053 53253
rect 28212 53201 28264 53253
rect 28423 53201 28475 53253
rect 28634 53201 28686 53253
rect 28845 53201 28897 53253
rect 29056 53201 29108 53253
rect 27790 51401 27842 51453
rect 28001 51401 28053 51453
rect 28212 51401 28264 51453
rect 28423 51401 28475 51453
rect 28634 51401 28686 51453
rect 28845 51401 28897 51453
rect 29056 51401 29108 51453
rect 27790 49601 27842 49653
rect 28001 49601 28053 49653
rect 28212 49601 28264 49653
rect 28423 49601 28475 49653
rect 28634 49601 28686 49653
rect 28845 49601 28897 49653
rect 29056 49601 29108 49653
rect 27790 47801 27842 47853
rect 28001 47801 28053 47853
rect 28212 47801 28264 47853
rect 28423 47801 28475 47853
rect 28634 47801 28686 47853
rect 28845 47801 28897 47853
rect 29056 47801 29108 47853
rect 27790 46001 27842 46053
rect 28001 46001 28053 46053
rect 28212 46001 28264 46053
rect 28423 46001 28475 46053
rect 28634 46001 28686 46053
rect 28845 46001 28897 46053
rect 29056 46001 29108 46053
rect 27790 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28686 44253
rect 28845 44201 28897 44253
rect 29056 44201 29108 44253
rect 27790 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28686 42453
rect 28845 42401 28897 42453
rect 29056 42401 29108 42453
rect 27790 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28686 40653
rect 28845 40601 28897 40653
rect 29056 40601 29108 40653
rect 27790 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28686 38853
rect 28845 38801 28897 38853
rect 29056 38801 29108 38853
rect 27790 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28686 37053
rect 28845 37001 28897 37053
rect 29056 37001 29108 37053
rect 56015 92801 56067 92853
rect 56226 92801 56278 92853
rect 56437 92801 56489 92853
rect 56648 92801 56700 92853
rect 56859 92801 56911 92853
rect 57070 92801 57122 92853
rect 57281 92801 57333 92853
rect 56015 91001 56067 91053
rect 56226 91001 56278 91053
rect 56437 91001 56489 91053
rect 56648 91001 56700 91053
rect 56859 91001 56911 91053
rect 57070 91001 57122 91053
rect 57281 91001 57333 91053
rect 56015 89201 56067 89253
rect 56226 89201 56278 89253
rect 56437 89201 56489 89253
rect 56648 89201 56700 89253
rect 56859 89201 56911 89253
rect 57070 89201 57122 89253
rect 57281 89201 57333 89253
rect 56015 87401 56067 87453
rect 56226 87401 56278 87453
rect 56437 87401 56489 87453
rect 56648 87401 56700 87453
rect 56859 87401 56911 87453
rect 57070 87401 57122 87453
rect 57281 87401 57333 87453
rect 56015 85601 56067 85653
rect 56226 85601 56278 85653
rect 56437 85601 56489 85653
rect 56648 85601 56700 85653
rect 56859 85601 56911 85653
rect 57070 85601 57122 85653
rect 57281 85601 57333 85653
rect 56015 83801 56067 83853
rect 56226 83801 56278 83853
rect 56437 83801 56489 83853
rect 56648 83801 56700 83853
rect 56859 83801 56911 83853
rect 57070 83801 57122 83853
rect 57281 83801 57333 83853
rect 56015 82001 56067 82053
rect 56226 82001 56278 82053
rect 56437 82001 56489 82053
rect 56648 82001 56700 82053
rect 56859 82001 56911 82053
rect 57070 82001 57122 82053
rect 57281 82001 57333 82053
rect 56015 80201 56067 80253
rect 56226 80201 56278 80253
rect 56437 80201 56489 80253
rect 56648 80201 56700 80253
rect 56859 80201 56911 80253
rect 57070 80201 57122 80253
rect 57281 80201 57333 80253
rect 56015 78401 56067 78453
rect 56226 78401 56278 78453
rect 56437 78401 56489 78453
rect 56648 78401 56700 78453
rect 56859 78401 56911 78453
rect 57070 78401 57122 78453
rect 57281 78401 57333 78453
rect 56015 76601 56067 76653
rect 56226 76601 56278 76653
rect 56437 76601 56489 76653
rect 56648 76601 56700 76653
rect 56859 76601 56911 76653
rect 57070 76601 57122 76653
rect 57281 76601 57333 76653
rect 56015 74801 56067 74853
rect 56226 74801 56278 74853
rect 56437 74801 56489 74853
rect 56648 74801 56700 74853
rect 56859 74801 56911 74853
rect 57070 74801 57122 74853
rect 57281 74801 57333 74853
rect 56015 73001 56067 73053
rect 56226 73001 56278 73053
rect 56437 73001 56489 73053
rect 56648 73001 56700 73053
rect 56859 73001 56911 73053
rect 57070 73001 57122 73053
rect 57281 73001 57333 73053
rect 56015 71201 56067 71253
rect 56226 71201 56278 71253
rect 56437 71201 56489 71253
rect 56648 71201 56700 71253
rect 56859 71201 56911 71253
rect 57070 71201 57122 71253
rect 57281 71201 57333 71253
rect 56015 69401 56067 69453
rect 56226 69401 56278 69453
rect 56437 69401 56489 69453
rect 56648 69401 56700 69453
rect 56859 69401 56911 69453
rect 57070 69401 57122 69453
rect 57281 69401 57333 69453
rect 56015 67601 56067 67653
rect 56226 67601 56278 67653
rect 56437 67601 56489 67653
rect 56648 67601 56700 67653
rect 56859 67601 56911 67653
rect 57070 67601 57122 67653
rect 57281 67601 57333 67653
rect 56015 65801 56067 65853
rect 56226 65801 56278 65853
rect 56437 65801 56489 65853
rect 56648 65801 56700 65853
rect 56859 65801 56911 65853
rect 57070 65801 57122 65853
rect 57281 65801 57333 65853
rect 56015 64001 56067 64053
rect 56226 64001 56278 64053
rect 56437 64001 56489 64053
rect 56648 64001 56700 64053
rect 56859 64001 56911 64053
rect 57070 64001 57122 64053
rect 57281 64001 57333 64053
rect 56015 62201 56067 62253
rect 56226 62201 56278 62253
rect 56437 62201 56489 62253
rect 56648 62201 56700 62253
rect 56859 62201 56911 62253
rect 57070 62201 57122 62253
rect 57281 62201 57333 62253
rect 56015 60401 56067 60453
rect 56226 60401 56278 60453
rect 56437 60401 56489 60453
rect 56648 60401 56700 60453
rect 56859 60401 56911 60453
rect 57070 60401 57122 60453
rect 57281 60401 57333 60453
rect 56015 58601 56067 58653
rect 56226 58601 56278 58653
rect 56437 58601 56489 58653
rect 56648 58601 56700 58653
rect 56859 58601 56911 58653
rect 57070 58601 57122 58653
rect 57281 58601 57333 58653
rect 56015 56801 56067 56853
rect 56226 56801 56278 56853
rect 56437 56801 56489 56853
rect 56648 56801 56700 56853
rect 56859 56801 56911 56853
rect 57070 56801 57122 56853
rect 57281 56801 57333 56853
rect 56015 55001 56067 55053
rect 56226 55001 56278 55053
rect 56437 55001 56489 55053
rect 56648 55001 56700 55053
rect 56859 55001 56911 55053
rect 57070 55001 57122 55053
rect 57281 55001 57333 55053
rect 56015 53201 56067 53253
rect 56226 53201 56278 53253
rect 56437 53201 56489 53253
rect 56648 53201 56700 53253
rect 56859 53201 56911 53253
rect 57070 53201 57122 53253
rect 57281 53201 57333 53253
rect 56015 51401 56067 51453
rect 56226 51401 56278 51453
rect 56437 51401 56489 51453
rect 56648 51401 56700 51453
rect 56859 51401 56911 51453
rect 57070 51401 57122 51453
rect 57281 51401 57333 51453
rect 56015 49601 56067 49653
rect 56226 49601 56278 49653
rect 56437 49601 56489 49653
rect 56648 49601 56700 49653
rect 56859 49601 56911 49653
rect 57070 49601 57122 49653
rect 57281 49601 57333 49653
rect 56015 47801 56067 47853
rect 56226 47801 56278 47853
rect 56437 47801 56489 47853
rect 56648 47801 56700 47853
rect 56859 47801 56911 47853
rect 57070 47801 57122 47853
rect 57281 47801 57333 47853
rect 56015 46001 56067 46053
rect 56226 46001 56278 46053
rect 56437 46001 56489 46053
rect 56648 46001 56700 46053
rect 56859 46001 56911 46053
rect 57070 46001 57122 46053
rect 57281 46001 57333 46053
rect 56015 44201 56067 44253
rect 56226 44201 56278 44253
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57333 44253
rect 56015 42401 56067 42453
rect 56226 42401 56278 42453
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57333 42453
rect 56015 40601 56067 40653
rect 56226 40601 56278 40653
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57333 40653
rect 56015 38801 56067 38853
rect 56226 38801 56278 38853
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57333 38853
rect 56015 37001 56067 37053
rect 56226 37001 56278 37053
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57333 37053
rect 60575 35338 60627 35494
rect 49908 6297 50064 6349
rect 51654 5147 51810 5199
rect 40623 3230 40779 3282
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 62150 1637 62306 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
<< metal2 >>
rect 282 96368 86090 96694
rect 706 95176 85666 96176
rect 706 282 1706 95176
rect 25313 26433 26039 94803
rect 26554 32126 26996 95176
rect 27387 94655 29146 94694
rect 27387 94599 27788 94655
rect 27844 94599 27999 94655
rect 28055 94599 28210 94655
rect 28266 94599 28421 94655
rect 28477 94599 28632 94655
rect 28688 94599 28843 94655
rect 28899 94599 29054 94655
rect 29110 94599 29146 94655
rect 27387 94560 29146 94599
rect 27387 92894 27828 94560
rect 29486 94485 30364 95176
rect 30769 94485 32888 95176
rect 35128 94485 36415 95176
rect 38953 94671 39618 95176
rect 48789 94485 49990 95176
rect 52226 94485 54354 95176
rect 54758 94485 55638 95176
rect 55977 94655 57371 94694
rect 55977 94599 56013 94655
rect 56069 94599 56224 94655
rect 56280 94599 56435 94655
rect 56491 94599 56646 94655
rect 56702 94599 56857 94655
rect 56913 94599 57068 94655
rect 57124 94599 57279 94655
rect 57335 94599 57371 94655
rect 55977 94560 57371 94599
rect 27387 92855 29146 92894
rect 27387 92799 27788 92855
rect 27844 92799 27999 92855
rect 28055 92799 28210 92855
rect 28266 92799 28421 92855
rect 28477 92799 28632 92855
rect 28688 92799 28843 92855
rect 28899 92799 29054 92855
rect 29110 92799 29146 92855
rect 27387 92760 29146 92799
rect 55977 92855 57371 92894
rect 55977 92799 56013 92855
rect 56069 92799 56224 92855
rect 56280 92799 56435 92855
rect 56491 92799 56646 92855
rect 56702 92799 56857 92855
rect 56913 92799 57068 92855
rect 57124 92799 57279 92855
rect 57335 92799 57371 92855
rect 55977 92760 57371 92799
rect 27387 91094 27828 92760
rect 27387 91055 29146 91094
rect 27387 90999 27788 91055
rect 27844 90999 27999 91055
rect 28055 90999 28210 91055
rect 28266 90999 28421 91055
rect 28477 90999 28632 91055
rect 28688 90999 28843 91055
rect 28899 90999 29054 91055
rect 29110 90999 29146 91055
rect 27387 90960 29146 90999
rect 55977 91055 57371 91094
rect 55977 90999 56013 91055
rect 56069 90999 56224 91055
rect 56280 90999 56435 91055
rect 56491 90999 56646 91055
rect 56702 90999 56857 91055
rect 56913 90999 57068 91055
rect 57124 90999 57279 91055
rect 57335 90999 57371 91055
rect 55977 90960 57371 90999
rect 27387 89294 27828 90960
rect 27387 89255 29146 89294
rect 27387 89199 27788 89255
rect 27844 89199 27999 89255
rect 28055 89199 28210 89255
rect 28266 89199 28421 89255
rect 28477 89199 28632 89255
rect 28688 89199 28843 89255
rect 28899 89199 29054 89255
rect 29110 89199 29146 89255
rect 27387 89160 29146 89199
rect 55977 89255 57371 89294
rect 55977 89199 56013 89255
rect 56069 89199 56224 89255
rect 56280 89199 56435 89255
rect 56491 89199 56646 89255
rect 56702 89199 56857 89255
rect 56913 89199 57068 89255
rect 57124 89199 57279 89255
rect 57335 89199 57371 89255
rect 55977 89160 57371 89199
rect 27387 87494 27828 89160
rect 27387 87455 29146 87494
rect 27387 87399 27788 87455
rect 27844 87399 27999 87455
rect 28055 87399 28210 87455
rect 28266 87399 28421 87455
rect 28477 87399 28632 87455
rect 28688 87399 28843 87455
rect 28899 87399 29054 87455
rect 29110 87399 29146 87455
rect 27387 87360 29146 87399
rect 55977 87455 57371 87494
rect 55977 87399 56013 87455
rect 56069 87399 56224 87455
rect 56280 87399 56435 87455
rect 56491 87399 56646 87455
rect 56702 87399 56857 87455
rect 56913 87399 57068 87455
rect 57124 87399 57279 87455
rect 57335 87399 57371 87455
rect 55977 87360 57371 87399
rect 27387 85694 27828 87360
rect 27387 85655 29146 85694
rect 27387 85599 27788 85655
rect 27844 85599 27999 85655
rect 28055 85599 28210 85655
rect 28266 85599 28421 85655
rect 28477 85599 28632 85655
rect 28688 85599 28843 85655
rect 28899 85599 29054 85655
rect 29110 85599 29146 85655
rect 27387 85560 29146 85599
rect 55977 85655 57371 85694
rect 55977 85599 56013 85655
rect 56069 85599 56224 85655
rect 56280 85599 56435 85655
rect 56491 85599 56646 85655
rect 56702 85599 56857 85655
rect 56913 85599 57068 85655
rect 57124 85599 57279 85655
rect 57335 85599 57371 85655
rect 55977 85560 57371 85599
rect 27387 83894 27828 85560
rect 27387 83855 29146 83894
rect 27387 83799 27788 83855
rect 27844 83799 27999 83855
rect 28055 83799 28210 83855
rect 28266 83799 28421 83855
rect 28477 83799 28632 83855
rect 28688 83799 28843 83855
rect 28899 83799 29054 83855
rect 29110 83799 29146 83855
rect 27387 83760 29146 83799
rect 55977 83855 57371 83894
rect 55977 83799 56013 83855
rect 56069 83799 56224 83855
rect 56280 83799 56435 83855
rect 56491 83799 56646 83855
rect 56702 83799 56857 83855
rect 56913 83799 57068 83855
rect 57124 83799 57279 83855
rect 57335 83799 57371 83855
rect 55977 83760 57371 83799
rect 27387 82094 27828 83760
rect 27387 82055 29146 82094
rect 27387 81999 27788 82055
rect 27844 81999 27999 82055
rect 28055 81999 28210 82055
rect 28266 81999 28421 82055
rect 28477 81999 28632 82055
rect 28688 81999 28843 82055
rect 28899 81999 29054 82055
rect 29110 81999 29146 82055
rect 27387 81960 29146 81999
rect 55977 82055 57371 82094
rect 55977 81999 56013 82055
rect 56069 81999 56224 82055
rect 56280 81999 56435 82055
rect 56491 81999 56646 82055
rect 56702 81999 56857 82055
rect 56913 81999 57068 82055
rect 57124 81999 57279 82055
rect 57335 81999 57371 82055
rect 55977 81960 57371 81999
rect 27387 80294 27828 81960
rect 27387 80255 29146 80294
rect 27387 80199 27788 80255
rect 27844 80199 27999 80255
rect 28055 80199 28210 80255
rect 28266 80199 28421 80255
rect 28477 80199 28632 80255
rect 28688 80199 28843 80255
rect 28899 80199 29054 80255
rect 29110 80199 29146 80255
rect 27387 80160 29146 80199
rect 55977 80255 57371 80294
rect 55977 80199 56013 80255
rect 56069 80199 56224 80255
rect 56280 80199 56435 80255
rect 56491 80199 56646 80255
rect 56702 80199 56857 80255
rect 56913 80199 57068 80255
rect 57124 80199 57279 80255
rect 57335 80199 57371 80255
rect 55977 80160 57371 80199
rect 27387 78494 27828 80160
rect 27387 78455 29146 78494
rect 27387 78399 27788 78455
rect 27844 78399 27999 78455
rect 28055 78399 28210 78455
rect 28266 78399 28421 78455
rect 28477 78399 28632 78455
rect 28688 78399 28843 78455
rect 28899 78399 29054 78455
rect 29110 78399 29146 78455
rect 27387 78360 29146 78399
rect 55977 78455 57371 78494
rect 55977 78399 56013 78455
rect 56069 78399 56224 78455
rect 56280 78399 56435 78455
rect 56491 78399 56646 78455
rect 56702 78399 56857 78455
rect 56913 78399 57068 78455
rect 57124 78399 57279 78455
rect 57335 78399 57371 78455
rect 55977 78360 57371 78399
rect 27387 76694 27828 78360
rect 27387 76655 29146 76694
rect 27387 76599 27788 76655
rect 27844 76599 27999 76655
rect 28055 76599 28210 76655
rect 28266 76599 28421 76655
rect 28477 76599 28632 76655
rect 28688 76599 28843 76655
rect 28899 76599 29054 76655
rect 29110 76599 29146 76655
rect 27387 76560 29146 76599
rect 55977 76655 57371 76694
rect 55977 76599 56013 76655
rect 56069 76599 56224 76655
rect 56280 76599 56435 76655
rect 56491 76599 56646 76655
rect 56702 76599 56857 76655
rect 56913 76599 57068 76655
rect 57124 76599 57279 76655
rect 57335 76599 57371 76655
rect 55977 76560 57371 76599
rect 27387 74894 27828 76560
rect 27387 74855 29146 74894
rect 27387 74799 27788 74855
rect 27844 74799 27999 74855
rect 28055 74799 28210 74855
rect 28266 74799 28421 74855
rect 28477 74799 28632 74855
rect 28688 74799 28843 74855
rect 28899 74799 29054 74855
rect 29110 74799 29146 74855
rect 27387 74760 29146 74799
rect 55977 74855 57371 74894
rect 55977 74799 56013 74855
rect 56069 74799 56224 74855
rect 56280 74799 56435 74855
rect 56491 74799 56646 74855
rect 56702 74799 56857 74855
rect 56913 74799 57068 74855
rect 57124 74799 57279 74855
rect 57335 74799 57371 74855
rect 55977 74760 57371 74799
rect 27387 73094 27828 74760
rect 27387 73055 29146 73094
rect 27387 72999 27788 73055
rect 27844 72999 27999 73055
rect 28055 72999 28210 73055
rect 28266 72999 28421 73055
rect 28477 72999 28632 73055
rect 28688 72999 28843 73055
rect 28899 72999 29054 73055
rect 29110 72999 29146 73055
rect 27387 72960 29146 72999
rect 55977 73055 57371 73094
rect 55977 72999 56013 73055
rect 56069 72999 56224 73055
rect 56280 72999 56435 73055
rect 56491 72999 56646 73055
rect 56702 72999 56857 73055
rect 56913 72999 57068 73055
rect 57124 72999 57279 73055
rect 57335 72999 57371 73055
rect 55977 72960 57371 72999
rect 27387 71294 27828 72960
rect 27387 71255 29146 71294
rect 27387 71199 27788 71255
rect 27844 71199 27999 71255
rect 28055 71199 28210 71255
rect 28266 71199 28421 71255
rect 28477 71199 28632 71255
rect 28688 71199 28843 71255
rect 28899 71199 29054 71255
rect 29110 71199 29146 71255
rect 27387 71160 29146 71199
rect 55977 71255 57371 71294
rect 55977 71199 56013 71255
rect 56069 71199 56224 71255
rect 56280 71199 56435 71255
rect 56491 71199 56646 71255
rect 56702 71199 56857 71255
rect 56913 71199 57068 71255
rect 57124 71199 57279 71255
rect 57335 71199 57371 71255
rect 55977 71160 57371 71199
rect 27387 69494 27828 71160
rect 27387 69455 29146 69494
rect 27387 69399 27788 69455
rect 27844 69399 27999 69455
rect 28055 69399 28210 69455
rect 28266 69399 28421 69455
rect 28477 69399 28632 69455
rect 28688 69399 28843 69455
rect 28899 69399 29054 69455
rect 29110 69399 29146 69455
rect 27387 69360 29146 69399
rect 55977 69455 57371 69494
rect 55977 69399 56013 69455
rect 56069 69399 56224 69455
rect 56280 69399 56435 69455
rect 56491 69399 56646 69455
rect 56702 69399 56857 69455
rect 56913 69399 57068 69455
rect 57124 69399 57279 69455
rect 57335 69399 57371 69455
rect 55977 69360 57371 69399
rect 27387 67694 27828 69360
rect 27387 67655 29146 67694
rect 27387 67599 27788 67655
rect 27844 67599 27999 67655
rect 28055 67599 28210 67655
rect 28266 67599 28421 67655
rect 28477 67599 28632 67655
rect 28688 67599 28843 67655
rect 28899 67599 29054 67655
rect 29110 67599 29146 67655
rect 27387 67560 29146 67599
rect 55977 67655 57371 67694
rect 55977 67599 56013 67655
rect 56069 67599 56224 67655
rect 56280 67599 56435 67655
rect 56491 67599 56646 67655
rect 56702 67599 56857 67655
rect 56913 67599 57068 67655
rect 57124 67599 57279 67655
rect 57335 67599 57371 67655
rect 55977 67560 57371 67599
rect 27387 65894 27828 67560
rect 27387 65855 29146 65894
rect 27387 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 29146 65855
rect 27387 65760 29146 65799
rect 55977 65855 57371 65894
rect 55977 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 57371 65855
rect 55977 65760 57371 65799
rect 27387 64094 27828 65760
rect 27387 64055 29146 64094
rect 27387 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 29146 64055
rect 27387 63960 29146 63999
rect 55977 64055 57371 64094
rect 55977 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 57371 64055
rect 55977 63960 57371 63999
rect 27387 62294 27828 63960
rect 27387 62255 29146 62294
rect 27387 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 29146 62255
rect 27387 62160 29146 62199
rect 55977 62255 57371 62294
rect 55977 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 57371 62255
rect 55977 62160 57371 62199
rect 27387 60494 27828 62160
rect 27387 60455 29146 60494
rect 27387 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 29146 60455
rect 27387 60360 29146 60399
rect 55977 60455 57371 60494
rect 55977 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 57371 60455
rect 55977 60360 57371 60399
rect 27387 58694 27828 60360
rect 27387 58655 29146 58694
rect 27387 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 29146 58655
rect 27387 58560 29146 58599
rect 55977 58655 57371 58694
rect 55977 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 57371 58655
rect 55977 58560 57371 58599
rect 27387 56894 27828 58560
rect 27387 56855 29146 56894
rect 27387 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 29146 56855
rect 27387 56760 29146 56799
rect 55977 56855 57371 56894
rect 55977 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 57371 56855
rect 55977 56760 57371 56799
rect 27387 55094 27828 56760
rect 27387 55055 29146 55094
rect 27387 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 29146 55055
rect 27387 54960 29146 54999
rect 55977 55055 57371 55094
rect 55977 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 57371 55055
rect 55977 54960 57371 54999
rect 27387 53294 27828 54960
rect 27387 53255 29146 53294
rect 27387 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 29146 53255
rect 27387 53160 29146 53199
rect 55977 53255 57371 53294
rect 55977 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 57371 53255
rect 55977 53160 57371 53199
rect 27387 51494 27828 53160
rect 27387 51455 29146 51494
rect 27387 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 29146 51455
rect 27387 51360 29146 51399
rect 55977 51455 57371 51494
rect 55977 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 57371 51455
rect 55977 51360 57371 51399
rect 27387 49694 27828 51360
rect 27387 49655 29146 49694
rect 27387 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 29146 49655
rect 27387 49560 29146 49599
rect 55977 49655 57371 49694
rect 55977 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 57371 49655
rect 55977 49560 57371 49599
rect 27387 47894 27828 49560
rect 27387 47855 29146 47894
rect 27387 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 29146 47855
rect 27387 47760 29146 47799
rect 55977 47855 57371 47894
rect 55977 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 57371 47855
rect 55977 47760 57371 47799
rect 27387 46094 27828 47760
rect 27387 46055 29146 46094
rect 27387 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 29146 46055
rect 27387 45960 29146 45999
rect 55977 46055 57371 46094
rect 55977 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 57371 46055
rect 55977 45960 57371 45999
rect 27387 44294 27828 45960
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 55977 44255 57371 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57371 44255
rect 55977 44160 57371 44199
rect 27387 42494 27828 44160
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 55977 42455 57371 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57371 42455
rect 55977 42360 57371 42399
rect 27387 40694 27828 42360
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 55977 40655 57371 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57371 40655
rect 55977 40560 57371 40599
rect 27387 38894 27828 40560
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 55977 38855 57371 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57371 38855
rect 55977 38760 57371 38799
rect 27387 37094 27828 38760
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 55977 37055 57371 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57371 37055
rect 55977 36960 57371 36999
rect 26554 32088 27163 32126
rect 26554 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27163 32088
rect 26554 31870 27163 32032
rect 26554 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27163 31870
rect 26554 31652 27163 31814
rect 26554 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27163 31652
rect 26554 31558 27163 31596
rect 26554 27382 26996 31558
rect 27387 26799 27828 36960
rect 36863 35881 37743 36650
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35761 41694 36096
rect 38596 35532 41694 35761
rect 38596 35516 38817 35532
rect 31615 35287 38817 35516
rect 41850 35425 42072 36096
rect 31615 33349 31836 35287
rect 39077 35197 42072 35425
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 36096
rect 31970 33349 32192 34943
rect 39755 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 36085
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 43205 34419
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 36085
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 43580 34083
rect 44646 35614 45735 35842
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 36096
rect 44997 35278 46112 35507
rect 46268 35681 46490 36096
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 36085
rect 47402 35171 47623 36096
rect 47779 35507 48001 36096
rect 48157 35842 48379 36096
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26581 27828 26743
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 27387 25028 27828 26525
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24810 27828 24972
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 26914 20570 27094 20580
rect 26914 20410 26924 20570
rect 27084 20410 27094 20570
rect 26914 20400 27094 20410
rect 26914 20226 27094 20236
rect 26914 20066 26924 20226
rect 27084 20066 27094 20226
rect 26914 20056 27094 20066
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 27387 7535 27828 24754
rect 57295 26799 57736 33519
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26581 57736 26743
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 49887 8953 50067 8963
rect 49887 8897 49897 8953
rect 50057 8897 50067 8953
rect 49887 8887 50067 8897
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6120 27828 7043
rect 49958 6361 50014 8887
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 5902 27828 6064
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 26823 5539 27163 5578
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5321 27163 5483
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3539 5001
rect 3445 1701 3539 4880
rect 11617 1701 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1701 12346 4684
rect 13538 1701 13594 4684
rect 14211 1701 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 23953 5135
rect 22345 4880 22621 5001
rect 22345 1701 22439 4880
rect 23859 3382 23953 5024
rect 26823 4528 27163 4567
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4310 27163 4472
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4215 27163 4254
rect 27387 3837 27828 5846
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3619 27828 3781
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 1701
rect 11533 0 11757 1701
rect 12206 0 12430 1701
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1701
rect 14127 0 14351 1701
rect 22279 0 22503 1701
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 3382
rect 27936 0 28160 3382
rect 29006 2524 29135 3418
rect 29247 3004 29377 3418
rect 29247 2768 29929 3004
rect 29006 0 29230 2524
rect 29705 0 29929 2768
rect 30859 0 31083 6229
rect 32552 0 32776 6229
rect 34243 0 34467 6229
rect 40588 3282 40812 3294
rect 40588 3230 40623 3282
rect 40779 3230 40812 3282
rect 40588 0 40812 3230
rect 43790 3050 43970 3060
rect 43790 2994 43800 3050
rect 43960 2994 43970 3050
rect 43790 2984 43970 2994
rect 50342 0 50566 7278
rect 51766 5211 51822 9801
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6120 57736 26525
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 5902 57736 6064
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 57295 3837 57736 5846
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 53772 3247 55669 3471
rect 53772 0 53996 3247
rect 55781 3024 55911 3418
rect 54417 2800 55911 3024
rect 54417 0 54641 2800
rect 56023 2540 56152 3418
rect 55164 2316 56152 2540
rect 55164 0 55388 2316
rect 56265 0 56489 3729
rect 57295 3619 57736 3781
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 32088 58351 95176
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31870 58351 32032
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31652 58351 31814
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 20570 58351 31596
rect 58791 26433 59517 94794
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 57909 20410 58048 20570
rect 58208 20410 58351 20570
rect 57909 20226 58351 20410
rect 57909 20066 58048 20226
rect 58208 20066 58351 20226
rect 57909 5539 58351 20066
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5321 58351 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 57909 4528 58351 5265
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4310 58351 4472
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 3524 58351 4254
rect 61447 5024 62085 5135
rect 71303 5073 71359 5140
rect 61447 0 61671 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 82103 5001 82197 5062
rect 82951 5024 83596 5135
rect 81921 4880 82197 5001
rect 81921 1701 82015 4880
rect 62115 1689 62339 1701
rect 62115 1637 62150 1689
rect 62306 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 5024
rect 84666 282 85666 95176
<< via2 >>
rect 27788 94653 27844 94655
rect 27788 94601 27790 94653
rect 27790 94601 27842 94653
rect 27842 94601 27844 94653
rect 27788 94599 27844 94601
rect 27999 94653 28055 94655
rect 27999 94601 28001 94653
rect 28001 94601 28053 94653
rect 28053 94601 28055 94653
rect 27999 94599 28055 94601
rect 28210 94653 28266 94655
rect 28210 94601 28212 94653
rect 28212 94601 28264 94653
rect 28264 94601 28266 94653
rect 28210 94599 28266 94601
rect 28421 94653 28477 94655
rect 28421 94601 28423 94653
rect 28423 94601 28475 94653
rect 28475 94601 28477 94653
rect 28421 94599 28477 94601
rect 28632 94653 28688 94655
rect 28632 94601 28634 94653
rect 28634 94601 28686 94653
rect 28686 94601 28688 94653
rect 28632 94599 28688 94601
rect 28843 94653 28899 94655
rect 28843 94601 28845 94653
rect 28845 94601 28897 94653
rect 28897 94601 28899 94653
rect 28843 94599 28899 94601
rect 29054 94653 29110 94655
rect 29054 94601 29056 94653
rect 29056 94601 29108 94653
rect 29108 94601 29110 94653
rect 29054 94599 29110 94601
rect 56013 94653 56069 94655
rect 56013 94601 56015 94653
rect 56015 94601 56067 94653
rect 56067 94601 56069 94653
rect 56013 94599 56069 94601
rect 56224 94653 56280 94655
rect 56224 94601 56226 94653
rect 56226 94601 56278 94653
rect 56278 94601 56280 94653
rect 56224 94599 56280 94601
rect 56435 94653 56491 94655
rect 56435 94601 56437 94653
rect 56437 94601 56489 94653
rect 56489 94601 56491 94653
rect 56435 94599 56491 94601
rect 56646 94653 56702 94655
rect 56646 94601 56648 94653
rect 56648 94601 56700 94653
rect 56700 94601 56702 94653
rect 56646 94599 56702 94601
rect 56857 94653 56913 94655
rect 56857 94601 56859 94653
rect 56859 94601 56911 94653
rect 56911 94601 56913 94653
rect 56857 94599 56913 94601
rect 57068 94653 57124 94655
rect 57068 94601 57070 94653
rect 57070 94601 57122 94653
rect 57122 94601 57124 94653
rect 57068 94599 57124 94601
rect 57279 94653 57335 94655
rect 57279 94601 57281 94653
rect 57281 94601 57333 94653
rect 57333 94601 57335 94653
rect 57279 94599 57335 94601
rect 27788 92853 27844 92855
rect 27788 92801 27790 92853
rect 27790 92801 27842 92853
rect 27842 92801 27844 92853
rect 27788 92799 27844 92801
rect 27999 92853 28055 92855
rect 27999 92801 28001 92853
rect 28001 92801 28053 92853
rect 28053 92801 28055 92853
rect 27999 92799 28055 92801
rect 28210 92853 28266 92855
rect 28210 92801 28212 92853
rect 28212 92801 28264 92853
rect 28264 92801 28266 92853
rect 28210 92799 28266 92801
rect 28421 92853 28477 92855
rect 28421 92801 28423 92853
rect 28423 92801 28475 92853
rect 28475 92801 28477 92853
rect 28421 92799 28477 92801
rect 28632 92853 28688 92855
rect 28632 92801 28634 92853
rect 28634 92801 28686 92853
rect 28686 92801 28688 92853
rect 28632 92799 28688 92801
rect 28843 92853 28899 92855
rect 28843 92801 28845 92853
rect 28845 92801 28897 92853
rect 28897 92801 28899 92853
rect 28843 92799 28899 92801
rect 29054 92853 29110 92855
rect 29054 92801 29056 92853
rect 29056 92801 29108 92853
rect 29108 92801 29110 92853
rect 29054 92799 29110 92801
rect 56013 92853 56069 92855
rect 56013 92801 56015 92853
rect 56015 92801 56067 92853
rect 56067 92801 56069 92853
rect 56013 92799 56069 92801
rect 56224 92853 56280 92855
rect 56224 92801 56226 92853
rect 56226 92801 56278 92853
rect 56278 92801 56280 92853
rect 56224 92799 56280 92801
rect 56435 92853 56491 92855
rect 56435 92801 56437 92853
rect 56437 92801 56489 92853
rect 56489 92801 56491 92853
rect 56435 92799 56491 92801
rect 56646 92853 56702 92855
rect 56646 92801 56648 92853
rect 56648 92801 56700 92853
rect 56700 92801 56702 92853
rect 56646 92799 56702 92801
rect 56857 92853 56913 92855
rect 56857 92801 56859 92853
rect 56859 92801 56911 92853
rect 56911 92801 56913 92853
rect 56857 92799 56913 92801
rect 57068 92853 57124 92855
rect 57068 92801 57070 92853
rect 57070 92801 57122 92853
rect 57122 92801 57124 92853
rect 57068 92799 57124 92801
rect 57279 92853 57335 92855
rect 57279 92801 57281 92853
rect 57281 92801 57333 92853
rect 57333 92801 57335 92853
rect 57279 92799 57335 92801
rect 27788 91053 27844 91055
rect 27788 91001 27790 91053
rect 27790 91001 27842 91053
rect 27842 91001 27844 91053
rect 27788 90999 27844 91001
rect 27999 91053 28055 91055
rect 27999 91001 28001 91053
rect 28001 91001 28053 91053
rect 28053 91001 28055 91053
rect 27999 90999 28055 91001
rect 28210 91053 28266 91055
rect 28210 91001 28212 91053
rect 28212 91001 28264 91053
rect 28264 91001 28266 91053
rect 28210 90999 28266 91001
rect 28421 91053 28477 91055
rect 28421 91001 28423 91053
rect 28423 91001 28475 91053
rect 28475 91001 28477 91053
rect 28421 90999 28477 91001
rect 28632 91053 28688 91055
rect 28632 91001 28634 91053
rect 28634 91001 28686 91053
rect 28686 91001 28688 91053
rect 28632 90999 28688 91001
rect 28843 91053 28899 91055
rect 28843 91001 28845 91053
rect 28845 91001 28897 91053
rect 28897 91001 28899 91053
rect 28843 90999 28899 91001
rect 29054 91053 29110 91055
rect 29054 91001 29056 91053
rect 29056 91001 29108 91053
rect 29108 91001 29110 91053
rect 29054 90999 29110 91001
rect 56013 91053 56069 91055
rect 56013 91001 56015 91053
rect 56015 91001 56067 91053
rect 56067 91001 56069 91053
rect 56013 90999 56069 91001
rect 56224 91053 56280 91055
rect 56224 91001 56226 91053
rect 56226 91001 56278 91053
rect 56278 91001 56280 91053
rect 56224 90999 56280 91001
rect 56435 91053 56491 91055
rect 56435 91001 56437 91053
rect 56437 91001 56489 91053
rect 56489 91001 56491 91053
rect 56435 90999 56491 91001
rect 56646 91053 56702 91055
rect 56646 91001 56648 91053
rect 56648 91001 56700 91053
rect 56700 91001 56702 91053
rect 56646 90999 56702 91001
rect 56857 91053 56913 91055
rect 56857 91001 56859 91053
rect 56859 91001 56911 91053
rect 56911 91001 56913 91053
rect 56857 90999 56913 91001
rect 57068 91053 57124 91055
rect 57068 91001 57070 91053
rect 57070 91001 57122 91053
rect 57122 91001 57124 91053
rect 57068 90999 57124 91001
rect 57279 91053 57335 91055
rect 57279 91001 57281 91053
rect 57281 91001 57333 91053
rect 57333 91001 57335 91053
rect 57279 90999 57335 91001
rect 27788 89253 27844 89255
rect 27788 89201 27790 89253
rect 27790 89201 27842 89253
rect 27842 89201 27844 89253
rect 27788 89199 27844 89201
rect 27999 89253 28055 89255
rect 27999 89201 28001 89253
rect 28001 89201 28053 89253
rect 28053 89201 28055 89253
rect 27999 89199 28055 89201
rect 28210 89253 28266 89255
rect 28210 89201 28212 89253
rect 28212 89201 28264 89253
rect 28264 89201 28266 89253
rect 28210 89199 28266 89201
rect 28421 89253 28477 89255
rect 28421 89201 28423 89253
rect 28423 89201 28475 89253
rect 28475 89201 28477 89253
rect 28421 89199 28477 89201
rect 28632 89253 28688 89255
rect 28632 89201 28634 89253
rect 28634 89201 28686 89253
rect 28686 89201 28688 89253
rect 28632 89199 28688 89201
rect 28843 89253 28899 89255
rect 28843 89201 28845 89253
rect 28845 89201 28897 89253
rect 28897 89201 28899 89253
rect 28843 89199 28899 89201
rect 29054 89253 29110 89255
rect 29054 89201 29056 89253
rect 29056 89201 29108 89253
rect 29108 89201 29110 89253
rect 29054 89199 29110 89201
rect 56013 89253 56069 89255
rect 56013 89201 56015 89253
rect 56015 89201 56067 89253
rect 56067 89201 56069 89253
rect 56013 89199 56069 89201
rect 56224 89253 56280 89255
rect 56224 89201 56226 89253
rect 56226 89201 56278 89253
rect 56278 89201 56280 89253
rect 56224 89199 56280 89201
rect 56435 89253 56491 89255
rect 56435 89201 56437 89253
rect 56437 89201 56489 89253
rect 56489 89201 56491 89253
rect 56435 89199 56491 89201
rect 56646 89253 56702 89255
rect 56646 89201 56648 89253
rect 56648 89201 56700 89253
rect 56700 89201 56702 89253
rect 56646 89199 56702 89201
rect 56857 89253 56913 89255
rect 56857 89201 56859 89253
rect 56859 89201 56911 89253
rect 56911 89201 56913 89253
rect 56857 89199 56913 89201
rect 57068 89253 57124 89255
rect 57068 89201 57070 89253
rect 57070 89201 57122 89253
rect 57122 89201 57124 89253
rect 57068 89199 57124 89201
rect 57279 89253 57335 89255
rect 57279 89201 57281 89253
rect 57281 89201 57333 89253
rect 57333 89201 57335 89253
rect 57279 89199 57335 89201
rect 27788 87453 27844 87455
rect 27788 87401 27790 87453
rect 27790 87401 27842 87453
rect 27842 87401 27844 87453
rect 27788 87399 27844 87401
rect 27999 87453 28055 87455
rect 27999 87401 28001 87453
rect 28001 87401 28053 87453
rect 28053 87401 28055 87453
rect 27999 87399 28055 87401
rect 28210 87453 28266 87455
rect 28210 87401 28212 87453
rect 28212 87401 28264 87453
rect 28264 87401 28266 87453
rect 28210 87399 28266 87401
rect 28421 87453 28477 87455
rect 28421 87401 28423 87453
rect 28423 87401 28475 87453
rect 28475 87401 28477 87453
rect 28421 87399 28477 87401
rect 28632 87453 28688 87455
rect 28632 87401 28634 87453
rect 28634 87401 28686 87453
rect 28686 87401 28688 87453
rect 28632 87399 28688 87401
rect 28843 87453 28899 87455
rect 28843 87401 28845 87453
rect 28845 87401 28897 87453
rect 28897 87401 28899 87453
rect 28843 87399 28899 87401
rect 29054 87453 29110 87455
rect 29054 87401 29056 87453
rect 29056 87401 29108 87453
rect 29108 87401 29110 87453
rect 29054 87399 29110 87401
rect 56013 87453 56069 87455
rect 56013 87401 56015 87453
rect 56015 87401 56067 87453
rect 56067 87401 56069 87453
rect 56013 87399 56069 87401
rect 56224 87453 56280 87455
rect 56224 87401 56226 87453
rect 56226 87401 56278 87453
rect 56278 87401 56280 87453
rect 56224 87399 56280 87401
rect 56435 87453 56491 87455
rect 56435 87401 56437 87453
rect 56437 87401 56489 87453
rect 56489 87401 56491 87453
rect 56435 87399 56491 87401
rect 56646 87453 56702 87455
rect 56646 87401 56648 87453
rect 56648 87401 56700 87453
rect 56700 87401 56702 87453
rect 56646 87399 56702 87401
rect 56857 87453 56913 87455
rect 56857 87401 56859 87453
rect 56859 87401 56911 87453
rect 56911 87401 56913 87453
rect 56857 87399 56913 87401
rect 57068 87453 57124 87455
rect 57068 87401 57070 87453
rect 57070 87401 57122 87453
rect 57122 87401 57124 87453
rect 57068 87399 57124 87401
rect 57279 87453 57335 87455
rect 57279 87401 57281 87453
rect 57281 87401 57333 87453
rect 57333 87401 57335 87453
rect 57279 87399 57335 87401
rect 27788 85653 27844 85655
rect 27788 85601 27790 85653
rect 27790 85601 27842 85653
rect 27842 85601 27844 85653
rect 27788 85599 27844 85601
rect 27999 85653 28055 85655
rect 27999 85601 28001 85653
rect 28001 85601 28053 85653
rect 28053 85601 28055 85653
rect 27999 85599 28055 85601
rect 28210 85653 28266 85655
rect 28210 85601 28212 85653
rect 28212 85601 28264 85653
rect 28264 85601 28266 85653
rect 28210 85599 28266 85601
rect 28421 85653 28477 85655
rect 28421 85601 28423 85653
rect 28423 85601 28475 85653
rect 28475 85601 28477 85653
rect 28421 85599 28477 85601
rect 28632 85653 28688 85655
rect 28632 85601 28634 85653
rect 28634 85601 28686 85653
rect 28686 85601 28688 85653
rect 28632 85599 28688 85601
rect 28843 85653 28899 85655
rect 28843 85601 28845 85653
rect 28845 85601 28897 85653
rect 28897 85601 28899 85653
rect 28843 85599 28899 85601
rect 29054 85653 29110 85655
rect 29054 85601 29056 85653
rect 29056 85601 29108 85653
rect 29108 85601 29110 85653
rect 29054 85599 29110 85601
rect 56013 85653 56069 85655
rect 56013 85601 56015 85653
rect 56015 85601 56067 85653
rect 56067 85601 56069 85653
rect 56013 85599 56069 85601
rect 56224 85653 56280 85655
rect 56224 85601 56226 85653
rect 56226 85601 56278 85653
rect 56278 85601 56280 85653
rect 56224 85599 56280 85601
rect 56435 85653 56491 85655
rect 56435 85601 56437 85653
rect 56437 85601 56489 85653
rect 56489 85601 56491 85653
rect 56435 85599 56491 85601
rect 56646 85653 56702 85655
rect 56646 85601 56648 85653
rect 56648 85601 56700 85653
rect 56700 85601 56702 85653
rect 56646 85599 56702 85601
rect 56857 85653 56913 85655
rect 56857 85601 56859 85653
rect 56859 85601 56911 85653
rect 56911 85601 56913 85653
rect 56857 85599 56913 85601
rect 57068 85653 57124 85655
rect 57068 85601 57070 85653
rect 57070 85601 57122 85653
rect 57122 85601 57124 85653
rect 57068 85599 57124 85601
rect 57279 85653 57335 85655
rect 57279 85601 57281 85653
rect 57281 85601 57333 85653
rect 57333 85601 57335 85653
rect 57279 85599 57335 85601
rect 27788 83853 27844 83855
rect 27788 83801 27790 83853
rect 27790 83801 27842 83853
rect 27842 83801 27844 83853
rect 27788 83799 27844 83801
rect 27999 83853 28055 83855
rect 27999 83801 28001 83853
rect 28001 83801 28053 83853
rect 28053 83801 28055 83853
rect 27999 83799 28055 83801
rect 28210 83853 28266 83855
rect 28210 83801 28212 83853
rect 28212 83801 28264 83853
rect 28264 83801 28266 83853
rect 28210 83799 28266 83801
rect 28421 83853 28477 83855
rect 28421 83801 28423 83853
rect 28423 83801 28475 83853
rect 28475 83801 28477 83853
rect 28421 83799 28477 83801
rect 28632 83853 28688 83855
rect 28632 83801 28634 83853
rect 28634 83801 28686 83853
rect 28686 83801 28688 83853
rect 28632 83799 28688 83801
rect 28843 83853 28899 83855
rect 28843 83801 28845 83853
rect 28845 83801 28897 83853
rect 28897 83801 28899 83853
rect 28843 83799 28899 83801
rect 29054 83853 29110 83855
rect 29054 83801 29056 83853
rect 29056 83801 29108 83853
rect 29108 83801 29110 83853
rect 29054 83799 29110 83801
rect 56013 83853 56069 83855
rect 56013 83801 56015 83853
rect 56015 83801 56067 83853
rect 56067 83801 56069 83853
rect 56013 83799 56069 83801
rect 56224 83853 56280 83855
rect 56224 83801 56226 83853
rect 56226 83801 56278 83853
rect 56278 83801 56280 83853
rect 56224 83799 56280 83801
rect 56435 83853 56491 83855
rect 56435 83801 56437 83853
rect 56437 83801 56489 83853
rect 56489 83801 56491 83853
rect 56435 83799 56491 83801
rect 56646 83853 56702 83855
rect 56646 83801 56648 83853
rect 56648 83801 56700 83853
rect 56700 83801 56702 83853
rect 56646 83799 56702 83801
rect 56857 83853 56913 83855
rect 56857 83801 56859 83853
rect 56859 83801 56911 83853
rect 56911 83801 56913 83853
rect 56857 83799 56913 83801
rect 57068 83853 57124 83855
rect 57068 83801 57070 83853
rect 57070 83801 57122 83853
rect 57122 83801 57124 83853
rect 57068 83799 57124 83801
rect 57279 83853 57335 83855
rect 57279 83801 57281 83853
rect 57281 83801 57333 83853
rect 57333 83801 57335 83853
rect 57279 83799 57335 83801
rect 27788 82053 27844 82055
rect 27788 82001 27790 82053
rect 27790 82001 27842 82053
rect 27842 82001 27844 82053
rect 27788 81999 27844 82001
rect 27999 82053 28055 82055
rect 27999 82001 28001 82053
rect 28001 82001 28053 82053
rect 28053 82001 28055 82053
rect 27999 81999 28055 82001
rect 28210 82053 28266 82055
rect 28210 82001 28212 82053
rect 28212 82001 28264 82053
rect 28264 82001 28266 82053
rect 28210 81999 28266 82001
rect 28421 82053 28477 82055
rect 28421 82001 28423 82053
rect 28423 82001 28475 82053
rect 28475 82001 28477 82053
rect 28421 81999 28477 82001
rect 28632 82053 28688 82055
rect 28632 82001 28634 82053
rect 28634 82001 28686 82053
rect 28686 82001 28688 82053
rect 28632 81999 28688 82001
rect 28843 82053 28899 82055
rect 28843 82001 28845 82053
rect 28845 82001 28897 82053
rect 28897 82001 28899 82053
rect 28843 81999 28899 82001
rect 29054 82053 29110 82055
rect 29054 82001 29056 82053
rect 29056 82001 29108 82053
rect 29108 82001 29110 82053
rect 29054 81999 29110 82001
rect 56013 82053 56069 82055
rect 56013 82001 56015 82053
rect 56015 82001 56067 82053
rect 56067 82001 56069 82053
rect 56013 81999 56069 82001
rect 56224 82053 56280 82055
rect 56224 82001 56226 82053
rect 56226 82001 56278 82053
rect 56278 82001 56280 82053
rect 56224 81999 56280 82001
rect 56435 82053 56491 82055
rect 56435 82001 56437 82053
rect 56437 82001 56489 82053
rect 56489 82001 56491 82053
rect 56435 81999 56491 82001
rect 56646 82053 56702 82055
rect 56646 82001 56648 82053
rect 56648 82001 56700 82053
rect 56700 82001 56702 82053
rect 56646 81999 56702 82001
rect 56857 82053 56913 82055
rect 56857 82001 56859 82053
rect 56859 82001 56911 82053
rect 56911 82001 56913 82053
rect 56857 81999 56913 82001
rect 57068 82053 57124 82055
rect 57068 82001 57070 82053
rect 57070 82001 57122 82053
rect 57122 82001 57124 82053
rect 57068 81999 57124 82001
rect 57279 82053 57335 82055
rect 57279 82001 57281 82053
rect 57281 82001 57333 82053
rect 57333 82001 57335 82053
rect 57279 81999 57335 82001
rect 27788 80253 27844 80255
rect 27788 80201 27790 80253
rect 27790 80201 27842 80253
rect 27842 80201 27844 80253
rect 27788 80199 27844 80201
rect 27999 80253 28055 80255
rect 27999 80201 28001 80253
rect 28001 80201 28053 80253
rect 28053 80201 28055 80253
rect 27999 80199 28055 80201
rect 28210 80253 28266 80255
rect 28210 80201 28212 80253
rect 28212 80201 28264 80253
rect 28264 80201 28266 80253
rect 28210 80199 28266 80201
rect 28421 80253 28477 80255
rect 28421 80201 28423 80253
rect 28423 80201 28475 80253
rect 28475 80201 28477 80253
rect 28421 80199 28477 80201
rect 28632 80253 28688 80255
rect 28632 80201 28634 80253
rect 28634 80201 28686 80253
rect 28686 80201 28688 80253
rect 28632 80199 28688 80201
rect 28843 80253 28899 80255
rect 28843 80201 28845 80253
rect 28845 80201 28897 80253
rect 28897 80201 28899 80253
rect 28843 80199 28899 80201
rect 29054 80253 29110 80255
rect 29054 80201 29056 80253
rect 29056 80201 29108 80253
rect 29108 80201 29110 80253
rect 29054 80199 29110 80201
rect 56013 80253 56069 80255
rect 56013 80201 56015 80253
rect 56015 80201 56067 80253
rect 56067 80201 56069 80253
rect 56013 80199 56069 80201
rect 56224 80253 56280 80255
rect 56224 80201 56226 80253
rect 56226 80201 56278 80253
rect 56278 80201 56280 80253
rect 56224 80199 56280 80201
rect 56435 80253 56491 80255
rect 56435 80201 56437 80253
rect 56437 80201 56489 80253
rect 56489 80201 56491 80253
rect 56435 80199 56491 80201
rect 56646 80253 56702 80255
rect 56646 80201 56648 80253
rect 56648 80201 56700 80253
rect 56700 80201 56702 80253
rect 56646 80199 56702 80201
rect 56857 80253 56913 80255
rect 56857 80201 56859 80253
rect 56859 80201 56911 80253
rect 56911 80201 56913 80253
rect 56857 80199 56913 80201
rect 57068 80253 57124 80255
rect 57068 80201 57070 80253
rect 57070 80201 57122 80253
rect 57122 80201 57124 80253
rect 57068 80199 57124 80201
rect 57279 80253 57335 80255
rect 57279 80201 57281 80253
rect 57281 80201 57333 80253
rect 57333 80201 57335 80253
rect 57279 80199 57335 80201
rect 27788 78453 27844 78455
rect 27788 78401 27790 78453
rect 27790 78401 27842 78453
rect 27842 78401 27844 78453
rect 27788 78399 27844 78401
rect 27999 78453 28055 78455
rect 27999 78401 28001 78453
rect 28001 78401 28053 78453
rect 28053 78401 28055 78453
rect 27999 78399 28055 78401
rect 28210 78453 28266 78455
rect 28210 78401 28212 78453
rect 28212 78401 28264 78453
rect 28264 78401 28266 78453
rect 28210 78399 28266 78401
rect 28421 78453 28477 78455
rect 28421 78401 28423 78453
rect 28423 78401 28475 78453
rect 28475 78401 28477 78453
rect 28421 78399 28477 78401
rect 28632 78453 28688 78455
rect 28632 78401 28634 78453
rect 28634 78401 28686 78453
rect 28686 78401 28688 78453
rect 28632 78399 28688 78401
rect 28843 78453 28899 78455
rect 28843 78401 28845 78453
rect 28845 78401 28897 78453
rect 28897 78401 28899 78453
rect 28843 78399 28899 78401
rect 29054 78453 29110 78455
rect 29054 78401 29056 78453
rect 29056 78401 29108 78453
rect 29108 78401 29110 78453
rect 29054 78399 29110 78401
rect 56013 78453 56069 78455
rect 56013 78401 56015 78453
rect 56015 78401 56067 78453
rect 56067 78401 56069 78453
rect 56013 78399 56069 78401
rect 56224 78453 56280 78455
rect 56224 78401 56226 78453
rect 56226 78401 56278 78453
rect 56278 78401 56280 78453
rect 56224 78399 56280 78401
rect 56435 78453 56491 78455
rect 56435 78401 56437 78453
rect 56437 78401 56489 78453
rect 56489 78401 56491 78453
rect 56435 78399 56491 78401
rect 56646 78453 56702 78455
rect 56646 78401 56648 78453
rect 56648 78401 56700 78453
rect 56700 78401 56702 78453
rect 56646 78399 56702 78401
rect 56857 78453 56913 78455
rect 56857 78401 56859 78453
rect 56859 78401 56911 78453
rect 56911 78401 56913 78453
rect 56857 78399 56913 78401
rect 57068 78453 57124 78455
rect 57068 78401 57070 78453
rect 57070 78401 57122 78453
rect 57122 78401 57124 78453
rect 57068 78399 57124 78401
rect 57279 78453 57335 78455
rect 57279 78401 57281 78453
rect 57281 78401 57333 78453
rect 57333 78401 57335 78453
rect 57279 78399 57335 78401
rect 27788 76653 27844 76655
rect 27788 76601 27790 76653
rect 27790 76601 27842 76653
rect 27842 76601 27844 76653
rect 27788 76599 27844 76601
rect 27999 76653 28055 76655
rect 27999 76601 28001 76653
rect 28001 76601 28053 76653
rect 28053 76601 28055 76653
rect 27999 76599 28055 76601
rect 28210 76653 28266 76655
rect 28210 76601 28212 76653
rect 28212 76601 28264 76653
rect 28264 76601 28266 76653
rect 28210 76599 28266 76601
rect 28421 76653 28477 76655
rect 28421 76601 28423 76653
rect 28423 76601 28475 76653
rect 28475 76601 28477 76653
rect 28421 76599 28477 76601
rect 28632 76653 28688 76655
rect 28632 76601 28634 76653
rect 28634 76601 28686 76653
rect 28686 76601 28688 76653
rect 28632 76599 28688 76601
rect 28843 76653 28899 76655
rect 28843 76601 28845 76653
rect 28845 76601 28897 76653
rect 28897 76601 28899 76653
rect 28843 76599 28899 76601
rect 29054 76653 29110 76655
rect 29054 76601 29056 76653
rect 29056 76601 29108 76653
rect 29108 76601 29110 76653
rect 29054 76599 29110 76601
rect 56013 76653 56069 76655
rect 56013 76601 56015 76653
rect 56015 76601 56067 76653
rect 56067 76601 56069 76653
rect 56013 76599 56069 76601
rect 56224 76653 56280 76655
rect 56224 76601 56226 76653
rect 56226 76601 56278 76653
rect 56278 76601 56280 76653
rect 56224 76599 56280 76601
rect 56435 76653 56491 76655
rect 56435 76601 56437 76653
rect 56437 76601 56489 76653
rect 56489 76601 56491 76653
rect 56435 76599 56491 76601
rect 56646 76653 56702 76655
rect 56646 76601 56648 76653
rect 56648 76601 56700 76653
rect 56700 76601 56702 76653
rect 56646 76599 56702 76601
rect 56857 76653 56913 76655
rect 56857 76601 56859 76653
rect 56859 76601 56911 76653
rect 56911 76601 56913 76653
rect 56857 76599 56913 76601
rect 57068 76653 57124 76655
rect 57068 76601 57070 76653
rect 57070 76601 57122 76653
rect 57122 76601 57124 76653
rect 57068 76599 57124 76601
rect 57279 76653 57335 76655
rect 57279 76601 57281 76653
rect 57281 76601 57333 76653
rect 57333 76601 57335 76653
rect 57279 76599 57335 76601
rect 27788 74853 27844 74855
rect 27788 74801 27790 74853
rect 27790 74801 27842 74853
rect 27842 74801 27844 74853
rect 27788 74799 27844 74801
rect 27999 74853 28055 74855
rect 27999 74801 28001 74853
rect 28001 74801 28053 74853
rect 28053 74801 28055 74853
rect 27999 74799 28055 74801
rect 28210 74853 28266 74855
rect 28210 74801 28212 74853
rect 28212 74801 28264 74853
rect 28264 74801 28266 74853
rect 28210 74799 28266 74801
rect 28421 74853 28477 74855
rect 28421 74801 28423 74853
rect 28423 74801 28475 74853
rect 28475 74801 28477 74853
rect 28421 74799 28477 74801
rect 28632 74853 28688 74855
rect 28632 74801 28634 74853
rect 28634 74801 28686 74853
rect 28686 74801 28688 74853
rect 28632 74799 28688 74801
rect 28843 74853 28899 74855
rect 28843 74801 28845 74853
rect 28845 74801 28897 74853
rect 28897 74801 28899 74853
rect 28843 74799 28899 74801
rect 29054 74853 29110 74855
rect 29054 74801 29056 74853
rect 29056 74801 29108 74853
rect 29108 74801 29110 74853
rect 29054 74799 29110 74801
rect 56013 74853 56069 74855
rect 56013 74801 56015 74853
rect 56015 74801 56067 74853
rect 56067 74801 56069 74853
rect 56013 74799 56069 74801
rect 56224 74853 56280 74855
rect 56224 74801 56226 74853
rect 56226 74801 56278 74853
rect 56278 74801 56280 74853
rect 56224 74799 56280 74801
rect 56435 74853 56491 74855
rect 56435 74801 56437 74853
rect 56437 74801 56489 74853
rect 56489 74801 56491 74853
rect 56435 74799 56491 74801
rect 56646 74853 56702 74855
rect 56646 74801 56648 74853
rect 56648 74801 56700 74853
rect 56700 74801 56702 74853
rect 56646 74799 56702 74801
rect 56857 74853 56913 74855
rect 56857 74801 56859 74853
rect 56859 74801 56911 74853
rect 56911 74801 56913 74853
rect 56857 74799 56913 74801
rect 57068 74853 57124 74855
rect 57068 74801 57070 74853
rect 57070 74801 57122 74853
rect 57122 74801 57124 74853
rect 57068 74799 57124 74801
rect 57279 74853 57335 74855
rect 57279 74801 57281 74853
rect 57281 74801 57333 74853
rect 57333 74801 57335 74853
rect 57279 74799 57335 74801
rect 27788 73053 27844 73055
rect 27788 73001 27790 73053
rect 27790 73001 27842 73053
rect 27842 73001 27844 73053
rect 27788 72999 27844 73001
rect 27999 73053 28055 73055
rect 27999 73001 28001 73053
rect 28001 73001 28053 73053
rect 28053 73001 28055 73053
rect 27999 72999 28055 73001
rect 28210 73053 28266 73055
rect 28210 73001 28212 73053
rect 28212 73001 28264 73053
rect 28264 73001 28266 73053
rect 28210 72999 28266 73001
rect 28421 73053 28477 73055
rect 28421 73001 28423 73053
rect 28423 73001 28475 73053
rect 28475 73001 28477 73053
rect 28421 72999 28477 73001
rect 28632 73053 28688 73055
rect 28632 73001 28634 73053
rect 28634 73001 28686 73053
rect 28686 73001 28688 73053
rect 28632 72999 28688 73001
rect 28843 73053 28899 73055
rect 28843 73001 28845 73053
rect 28845 73001 28897 73053
rect 28897 73001 28899 73053
rect 28843 72999 28899 73001
rect 29054 73053 29110 73055
rect 29054 73001 29056 73053
rect 29056 73001 29108 73053
rect 29108 73001 29110 73053
rect 29054 72999 29110 73001
rect 56013 73053 56069 73055
rect 56013 73001 56015 73053
rect 56015 73001 56067 73053
rect 56067 73001 56069 73053
rect 56013 72999 56069 73001
rect 56224 73053 56280 73055
rect 56224 73001 56226 73053
rect 56226 73001 56278 73053
rect 56278 73001 56280 73053
rect 56224 72999 56280 73001
rect 56435 73053 56491 73055
rect 56435 73001 56437 73053
rect 56437 73001 56489 73053
rect 56489 73001 56491 73053
rect 56435 72999 56491 73001
rect 56646 73053 56702 73055
rect 56646 73001 56648 73053
rect 56648 73001 56700 73053
rect 56700 73001 56702 73053
rect 56646 72999 56702 73001
rect 56857 73053 56913 73055
rect 56857 73001 56859 73053
rect 56859 73001 56911 73053
rect 56911 73001 56913 73053
rect 56857 72999 56913 73001
rect 57068 73053 57124 73055
rect 57068 73001 57070 73053
rect 57070 73001 57122 73053
rect 57122 73001 57124 73053
rect 57068 72999 57124 73001
rect 57279 73053 57335 73055
rect 57279 73001 57281 73053
rect 57281 73001 57333 73053
rect 57333 73001 57335 73053
rect 57279 72999 57335 73001
rect 27788 71253 27844 71255
rect 27788 71201 27790 71253
rect 27790 71201 27842 71253
rect 27842 71201 27844 71253
rect 27788 71199 27844 71201
rect 27999 71253 28055 71255
rect 27999 71201 28001 71253
rect 28001 71201 28053 71253
rect 28053 71201 28055 71253
rect 27999 71199 28055 71201
rect 28210 71253 28266 71255
rect 28210 71201 28212 71253
rect 28212 71201 28264 71253
rect 28264 71201 28266 71253
rect 28210 71199 28266 71201
rect 28421 71253 28477 71255
rect 28421 71201 28423 71253
rect 28423 71201 28475 71253
rect 28475 71201 28477 71253
rect 28421 71199 28477 71201
rect 28632 71253 28688 71255
rect 28632 71201 28634 71253
rect 28634 71201 28686 71253
rect 28686 71201 28688 71253
rect 28632 71199 28688 71201
rect 28843 71253 28899 71255
rect 28843 71201 28845 71253
rect 28845 71201 28897 71253
rect 28897 71201 28899 71253
rect 28843 71199 28899 71201
rect 29054 71253 29110 71255
rect 29054 71201 29056 71253
rect 29056 71201 29108 71253
rect 29108 71201 29110 71253
rect 29054 71199 29110 71201
rect 56013 71253 56069 71255
rect 56013 71201 56015 71253
rect 56015 71201 56067 71253
rect 56067 71201 56069 71253
rect 56013 71199 56069 71201
rect 56224 71253 56280 71255
rect 56224 71201 56226 71253
rect 56226 71201 56278 71253
rect 56278 71201 56280 71253
rect 56224 71199 56280 71201
rect 56435 71253 56491 71255
rect 56435 71201 56437 71253
rect 56437 71201 56489 71253
rect 56489 71201 56491 71253
rect 56435 71199 56491 71201
rect 56646 71253 56702 71255
rect 56646 71201 56648 71253
rect 56648 71201 56700 71253
rect 56700 71201 56702 71253
rect 56646 71199 56702 71201
rect 56857 71253 56913 71255
rect 56857 71201 56859 71253
rect 56859 71201 56911 71253
rect 56911 71201 56913 71253
rect 56857 71199 56913 71201
rect 57068 71253 57124 71255
rect 57068 71201 57070 71253
rect 57070 71201 57122 71253
rect 57122 71201 57124 71253
rect 57068 71199 57124 71201
rect 57279 71253 57335 71255
rect 57279 71201 57281 71253
rect 57281 71201 57333 71253
rect 57333 71201 57335 71253
rect 57279 71199 57335 71201
rect 27788 69453 27844 69455
rect 27788 69401 27790 69453
rect 27790 69401 27842 69453
rect 27842 69401 27844 69453
rect 27788 69399 27844 69401
rect 27999 69453 28055 69455
rect 27999 69401 28001 69453
rect 28001 69401 28053 69453
rect 28053 69401 28055 69453
rect 27999 69399 28055 69401
rect 28210 69453 28266 69455
rect 28210 69401 28212 69453
rect 28212 69401 28264 69453
rect 28264 69401 28266 69453
rect 28210 69399 28266 69401
rect 28421 69453 28477 69455
rect 28421 69401 28423 69453
rect 28423 69401 28475 69453
rect 28475 69401 28477 69453
rect 28421 69399 28477 69401
rect 28632 69453 28688 69455
rect 28632 69401 28634 69453
rect 28634 69401 28686 69453
rect 28686 69401 28688 69453
rect 28632 69399 28688 69401
rect 28843 69453 28899 69455
rect 28843 69401 28845 69453
rect 28845 69401 28897 69453
rect 28897 69401 28899 69453
rect 28843 69399 28899 69401
rect 29054 69453 29110 69455
rect 29054 69401 29056 69453
rect 29056 69401 29108 69453
rect 29108 69401 29110 69453
rect 29054 69399 29110 69401
rect 56013 69453 56069 69455
rect 56013 69401 56015 69453
rect 56015 69401 56067 69453
rect 56067 69401 56069 69453
rect 56013 69399 56069 69401
rect 56224 69453 56280 69455
rect 56224 69401 56226 69453
rect 56226 69401 56278 69453
rect 56278 69401 56280 69453
rect 56224 69399 56280 69401
rect 56435 69453 56491 69455
rect 56435 69401 56437 69453
rect 56437 69401 56489 69453
rect 56489 69401 56491 69453
rect 56435 69399 56491 69401
rect 56646 69453 56702 69455
rect 56646 69401 56648 69453
rect 56648 69401 56700 69453
rect 56700 69401 56702 69453
rect 56646 69399 56702 69401
rect 56857 69453 56913 69455
rect 56857 69401 56859 69453
rect 56859 69401 56911 69453
rect 56911 69401 56913 69453
rect 56857 69399 56913 69401
rect 57068 69453 57124 69455
rect 57068 69401 57070 69453
rect 57070 69401 57122 69453
rect 57122 69401 57124 69453
rect 57068 69399 57124 69401
rect 57279 69453 57335 69455
rect 57279 69401 57281 69453
rect 57281 69401 57333 69453
rect 57333 69401 57335 69453
rect 57279 69399 57335 69401
rect 27788 67653 27844 67655
rect 27788 67601 27790 67653
rect 27790 67601 27842 67653
rect 27842 67601 27844 67653
rect 27788 67599 27844 67601
rect 27999 67653 28055 67655
rect 27999 67601 28001 67653
rect 28001 67601 28053 67653
rect 28053 67601 28055 67653
rect 27999 67599 28055 67601
rect 28210 67653 28266 67655
rect 28210 67601 28212 67653
rect 28212 67601 28264 67653
rect 28264 67601 28266 67653
rect 28210 67599 28266 67601
rect 28421 67653 28477 67655
rect 28421 67601 28423 67653
rect 28423 67601 28475 67653
rect 28475 67601 28477 67653
rect 28421 67599 28477 67601
rect 28632 67653 28688 67655
rect 28632 67601 28634 67653
rect 28634 67601 28686 67653
rect 28686 67601 28688 67653
rect 28632 67599 28688 67601
rect 28843 67653 28899 67655
rect 28843 67601 28845 67653
rect 28845 67601 28897 67653
rect 28897 67601 28899 67653
rect 28843 67599 28899 67601
rect 29054 67653 29110 67655
rect 29054 67601 29056 67653
rect 29056 67601 29108 67653
rect 29108 67601 29110 67653
rect 29054 67599 29110 67601
rect 56013 67653 56069 67655
rect 56013 67601 56015 67653
rect 56015 67601 56067 67653
rect 56067 67601 56069 67653
rect 56013 67599 56069 67601
rect 56224 67653 56280 67655
rect 56224 67601 56226 67653
rect 56226 67601 56278 67653
rect 56278 67601 56280 67653
rect 56224 67599 56280 67601
rect 56435 67653 56491 67655
rect 56435 67601 56437 67653
rect 56437 67601 56489 67653
rect 56489 67601 56491 67653
rect 56435 67599 56491 67601
rect 56646 67653 56702 67655
rect 56646 67601 56648 67653
rect 56648 67601 56700 67653
rect 56700 67601 56702 67653
rect 56646 67599 56702 67601
rect 56857 67653 56913 67655
rect 56857 67601 56859 67653
rect 56859 67601 56911 67653
rect 56911 67601 56913 67653
rect 56857 67599 56913 67601
rect 57068 67653 57124 67655
rect 57068 67601 57070 67653
rect 57070 67601 57122 67653
rect 57122 67601 57124 67653
rect 57068 67599 57124 67601
rect 57279 67653 57335 67655
rect 57279 67601 57281 67653
rect 57281 67601 57333 67653
rect 57333 67601 57335 67653
rect 57279 67599 57335 67601
rect 27788 65853 27844 65855
rect 27788 65801 27790 65853
rect 27790 65801 27842 65853
rect 27842 65801 27844 65853
rect 27788 65799 27844 65801
rect 27999 65853 28055 65855
rect 27999 65801 28001 65853
rect 28001 65801 28053 65853
rect 28053 65801 28055 65853
rect 27999 65799 28055 65801
rect 28210 65853 28266 65855
rect 28210 65801 28212 65853
rect 28212 65801 28264 65853
rect 28264 65801 28266 65853
rect 28210 65799 28266 65801
rect 28421 65853 28477 65855
rect 28421 65801 28423 65853
rect 28423 65801 28475 65853
rect 28475 65801 28477 65853
rect 28421 65799 28477 65801
rect 28632 65853 28688 65855
rect 28632 65801 28634 65853
rect 28634 65801 28686 65853
rect 28686 65801 28688 65853
rect 28632 65799 28688 65801
rect 28843 65853 28899 65855
rect 28843 65801 28845 65853
rect 28845 65801 28897 65853
rect 28897 65801 28899 65853
rect 28843 65799 28899 65801
rect 29054 65853 29110 65855
rect 29054 65801 29056 65853
rect 29056 65801 29108 65853
rect 29108 65801 29110 65853
rect 29054 65799 29110 65801
rect 56013 65853 56069 65855
rect 56013 65801 56015 65853
rect 56015 65801 56067 65853
rect 56067 65801 56069 65853
rect 56013 65799 56069 65801
rect 56224 65853 56280 65855
rect 56224 65801 56226 65853
rect 56226 65801 56278 65853
rect 56278 65801 56280 65853
rect 56224 65799 56280 65801
rect 56435 65853 56491 65855
rect 56435 65801 56437 65853
rect 56437 65801 56489 65853
rect 56489 65801 56491 65853
rect 56435 65799 56491 65801
rect 56646 65853 56702 65855
rect 56646 65801 56648 65853
rect 56648 65801 56700 65853
rect 56700 65801 56702 65853
rect 56646 65799 56702 65801
rect 56857 65853 56913 65855
rect 56857 65801 56859 65853
rect 56859 65801 56911 65853
rect 56911 65801 56913 65853
rect 56857 65799 56913 65801
rect 57068 65853 57124 65855
rect 57068 65801 57070 65853
rect 57070 65801 57122 65853
rect 57122 65801 57124 65853
rect 57068 65799 57124 65801
rect 57279 65853 57335 65855
rect 57279 65801 57281 65853
rect 57281 65801 57333 65853
rect 57333 65801 57335 65853
rect 57279 65799 57335 65801
rect 27788 64053 27844 64055
rect 27788 64001 27790 64053
rect 27790 64001 27842 64053
rect 27842 64001 27844 64053
rect 27788 63999 27844 64001
rect 27999 64053 28055 64055
rect 27999 64001 28001 64053
rect 28001 64001 28053 64053
rect 28053 64001 28055 64053
rect 27999 63999 28055 64001
rect 28210 64053 28266 64055
rect 28210 64001 28212 64053
rect 28212 64001 28264 64053
rect 28264 64001 28266 64053
rect 28210 63999 28266 64001
rect 28421 64053 28477 64055
rect 28421 64001 28423 64053
rect 28423 64001 28475 64053
rect 28475 64001 28477 64053
rect 28421 63999 28477 64001
rect 28632 64053 28688 64055
rect 28632 64001 28634 64053
rect 28634 64001 28686 64053
rect 28686 64001 28688 64053
rect 28632 63999 28688 64001
rect 28843 64053 28899 64055
rect 28843 64001 28845 64053
rect 28845 64001 28897 64053
rect 28897 64001 28899 64053
rect 28843 63999 28899 64001
rect 29054 64053 29110 64055
rect 29054 64001 29056 64053
rect 29056 64001 29108 64053
rect 29108 64001 29110 64053
rect 29054 63999 29110 64001
rect 56013 64053 56069 64055
rect 56013 64001 56015 64053
rect 56015 64001 56067 64053
rect 56067 64001 56069 64053
rect 56013 63999 56069 64001
rect 56224 64053 56280 64055
rect 56224 64001 56226 64053
rect 56226 64001 56278 64053
rect 56278 64001 56280 64053
rect 56224 63999 56280 64001
rect 56435 64053 56491 64055
rect 56435 64001 56437 64053
rect 56437 64001 56489 64053
rect 56489 64001 56491 64053
rect 56435 63999 56491 64001
rect 56646 64053 56702 64055
rect 56646 64001 56648 64053
rect 56648 64001 56700 64053
rect 56700 64001 56702 64053
rect 56646 63999 56702 64001
rect 56857 64053 56913 64055
rect 56857 64001 56859 64053
rect 56859 64001 56911 64053
rect 56911 64001 56913 64053
rect 56857 63999 56913 64001
rect 57068 64053 57124 64055
rect 57068 64001 57070 64053
rect 57070 64001 57122 64053
rect 57122 64001 57124 64053
rect 57068 63999 57124 64001
rect 57279 64053 57335 64055
rect 57279 64001 57281 64053
rect 57281 64001 57333 64053
rect 57333 64001 57335 64053
rect 57279 63999 57335 64001
rect 27788 62253 27844 62255
rect 27788 62201 27790 62253
rect 27790 62201 27842 62253
rect 27842 62201 27844 62253
rect 27788 62199 27844 62201
rect 27999 62253 28055 62255
rect 27999 62201 28001 62253
rect 28001 62201 28053 62253
rect 28053 62201 28055 62253
rect 27999 62199 28055 62201
rect 28210 62253 28266 62255
rect 28210 62201 28212 62253
rect 28212 62201 28264 62253
rect 28264 62201 28266 62253
rect 28210 62199 28266 62201
rect 28421 62253 28477 62255
rect 28421 62201 28423 62253
rect 28423 62201 28475 62253
rect 28475 62201 28477 62253
rect 28421 62199 28477 62201
rect 28632 62253 28688 62255
rect 28632 62201 28634 62253
rect 28634 62201 28686 62253
rect 28686 62201 28688 62253
rect 28632 62199 28688 62201
rect 28843 62253 28899 62255
rect 28843 62201 28845 62253
rect 28845 62201 28897 62253
rect 28897 62201 28899 62253
rect 28843 62199 28899 62201
rect 29054 62253 29110 62255
rect 29054 62201 29056 62253
rect 29056 62201 29108 62253
rect 29108 62201 29110 62253
rect 29054 62199 29110 62201
rect 56013 62253 56069 62255
rect 56013 62201 56015 62253
rect 56015 62201 56067 62253
rect 56067 62201 56069 62253
rect 56013 62199 56069 62201
rect 56224 62253 56280 62255
rect 56224 62201 56226 62253
rect 56226 62201 56278 62253
rect 56278 62201 56280 62253
rect 56224 62199 56280 62201
rect 56435 62253 56491 62255
rect 56435 62201 56437 62253
rect 56437 62201 56489 62253
rect 56489 62201 56491 62253
rect 56435 62199 56491 62201
rect 56646 62253 56702 62255
rect 56646 62201 56648 62253
rect 56648 62201 56700 62253
rect 56700 62201 56702 62253
rect 56646 62199 56702 62201
rect 56857 62253 56913 62255
rect 56857 62201 56859 62253
rect 56859 62201 56911 62253
rect 56911 62201 56913 62253
rect 56857 62199 56913 62201
rect 57068 62253 57124 62255
rect 57068 62201 57070 62253
rect 57070 62201 57122 62253
rect 57122 62201 57124 62253
rect 57068 62199 57124 62201
rect 57279 62253 57335 62255
rect 57279 62201 57281 62253
rect 57281 62201 57333 62253
rect 57333 62201 57335 62253
rect 57279 62199 57335 62201
rect 27788 60453 27844 60455
rect 27788 60401 27790 60453
rect 27790 60401 27842 60453
rect 27842 60401 27844 60453
rect 27788 60399 27844 60401
rect 27999 60453 28055 60455
rect 27999 60401 28001 60453
rect 28001 60401 28053 60453
rect 28053 60401 28055 60453
rect 27999 60399 28055 60401
rect 28210 60453 28266 60455
rect 28210 60401 28212 60453
rect 28212 60401 28264 60453
rect 28264 60401 28266 60453
rect 28210 60399 28266 60401
rect 28421 60453 28477 60455
rect 28421 60401 28423 60453
rect 28423 60401 28475 60453
rect 28475 60401 28477 60453
rect 28421 60399 28477 60401
rect 28632 60453 28688 60455
rect 28632 60401 28634 60453
rect 28634 60401 28686 60453
rect 28686 60401 28688 60453
rect 28632 60399 28688 60401
rect 28843 60453 28899 60455
rect 28843 60401 28845 60453
rect 28845 60401 28897 60453
rect 28897 60401 28899 60453
rect 28843 60399 28899 60401
rect 29054 60453 29110 60455
rect 29054 60401 29056 60453
rect 29056 60401 29108 60453
rect 29108 60401 29110 60453
rect 29054 60399 29110 60401
rect 56013 60453 56069 60455
rect 56013 60401 56015 60453
rect 56015 60401 56067 60453
rect 56067 60401 56069 60453
rect 56013 60399 56069 60401
rect 56224 60453 56280 60455
rect 56224 60401 56226 60453
rect 56226 60401 56278 60453
rect 56278 60401 56280 60453
rect 56224 60399 56280 60401
rect 56435 60453 56491 60455
rect 56435 60401 56437 60453
rect 56437 60401 56489 60453
rect 56489 60401 56491 60453
rect 56435 60399 56491 60401
rect 56646 60453 56702 60455
rect 56646 60401 56648 60453
rect 56648 60401 56700 60453
rect 56700 60401 56702 60453
rect 56646 60399 56702 60401
rect 56857 60453 56913 60455
rect 56857 60401 56859 60453
rect 56859 60401 56911 60453
rect 56911 60401 56913 60453
rect 56857 60399 56913 60401
rect 57068 60453 57124 60455
rect 57068 60401 57070 60453
rect 57070 60401 57122 60453
rect 57122 60401 57124 60453
rect 57068 60399 57124 60401
rect 57279 60453 57335 60455
rect 57279 60401 57281 60453
rect 57281 60401 57333 60453
rect 57333 60401 57335 60453
rect 57279 60399 57335 60401
rect 27788 58653 27844 58655
rect 27788 58601 27790 58653
rect 27790 58601 27842 58653
rect 27842 58601 27844 58653
rect 27788 58599 27844 58601
rect 27999 58653 28055 58655
rect 27999 58601 28001 58653
rect 28001 58601 28053 58653
rect 28053 58601 28055 58653
rect 27999 58599 28055 58601
rect 28210 58653 28266 58655
rect 28210 58601 28212 58653
rect 28212 58601 28264 58653
rect 28264 58601 28266 58653
rect 28210 58599 28266 58601
rect 28421 58653 28477 58655
rect 28421 58601 28423 58653
rect 28423 58601 28475 58653
rect 28475 58601 28477 58653
rect 28421 58599 28477 58601
rect 28632 58653 28688 58655
rect 28632 58601 28634 58653
rect 28634 58601 28686 58653
rect 28686 58601 28688 58653
rect 28632 58599 28688 58601
rect 28843 58653 28899 58655
rect 28843 58601 28845 58653
rect 28845 58601 28897 58653
rect 28897 58601 28899 58653
rect 28843 58599 28899 58601
rect 29054 58653 29110 58655
rect 29054 58601 29056 58653
rect 29056 58601 29108 58653
rect 29108 58601 29110 58653
rect 29054 58599 29110 58601
rect 56013 58653 56069 58655
rect 56013 58601 56015 58653
rect 56015 58601 56067 58653
rect 56067 58601 56069 58653
rect 56013 58599 56069 58601
rect 56224 58653 56280 58655
rect 56224 58601 56226 58653
rect 56226 58601 56278 58653
rect 56278 58601 56280 58653
rect 56224 58599 56280 58601
rect 56435 58653 56491 58655
rect 56435 58601 56437 58653
rect 56437 58601 56489 58653
rect 56489 58601 56491 58653
rect 56435 58599 56491 58601
rect 56646 58653 56702 58655
rect 56646 58601 56648 58653
rect 56648 58601 56700 58653
rect 56700 58601 56702 58653
rect 56646 58599 56702 58601
rect 56857 58653 56913 58655
rect 56857 58601 56859 58653
rect 56859 58601 56911 58653
rect 56911 58601 56913 58653
rect 56857 58599 56913 58601
rect 57068 58653 57124 58655
rect 57068 58601 57070 58653
rect 57070 58601 57122 58653
rect 57122 58601 57124 58653
rect 57068 58599 57124 58601
rect 57279 58653 57335 58655
rect 57279 58601 57281 58653
rect 57281 58601 57333 58653
rect 57333 58601 57335 58653
rect 57279 58599 57335 58601
rect 27788 56853 27844 56855
rect 27788 56801 27790 56853
rect 27790 56801 27842 56853
rect 27842 56801 27844 56853
rect 27788 56799 27844 56801
rect 27999 56853 28055 56855
rect 27999 56801 28001 56853
rect 28001 56801 28053 56853
rect 28053 56801 28055 56853
rect 27999 56799 28055 56801
rect 28210 56853 28266 56855
rect 28210 56801 28212 56853
rect 28212 56801 28264 56853
rect 28264 56801 28266 56853
rect 28210 56799 28266 56801
rect 28421 56853 28477 56855
rect 28421 56801 28423 56853
rect 28423 56801 28475 56853
rect 28475 56801 28477 56853
rect 28421 56799 28477 56801
rect 28632 56853 28688 56855
rect 28632 56801 28634 56853
rect 28634 56801 28686 56853
rect 28686 56801 28688 56853
rect 28632 56799 28688 56801
rect 28843 56853 28899 56855
rect 28843 56801 28845 56853
rect 28845 56801 28897 56853
rect 28897 56801 28899 56853
rect 28843 56799 28899 56801
rect 29054 56853 29110 56855
rect 29054 56801 29056 56853
rect 29056 56801 29108 56853
rect 29108 56801 29110 56853
rect 29054 56799 29110 56801
rect 56013 56853 56069 56855
rect 56013 56801 56015 56853
rect 56015 56801 56067 56853
rect 56067 56801 56069 56853
rect 56013 56799 56069 56801
rect 56224 56853 56280 56855
rect 56224 56801 56226 56853
rect 56226 56801 56278 56853
rect 56278 56801 56280 56853
rect 56224 56799 56280 56801
rect 56435 56853 56491 56855
rect 56435 56801 56437 56853
rect 56437 56801 56489 56853
rect 56489 56801 56491 56853
rect 56435 56799 56491 56801
rect 56646 56853 56702 56855
rect 56646 56801 56648 56853
rect 56648 56801 56700 56853
rect 56700 56801 56702 56853
rect 56646 56799 56702 56801
rect 56857 56853 56913 56855
rect 56857 56801 56859 56853
rect 56859 56801 56911 56853
rect 56911 56801 56913 56853
rect 56857 56799 56913 56801
rect 57068 56853 57124 56855
rect 57068 56801 57070 56853
rect 57070 56801 57122 56853
rect 57122 56801 57124 56853
rect 57068 56799 57124 56801
rect 57279 56853 57335 56855
rect 57279 56801 57281 56853
rect 57281 56801 57333 56853
rect 57333 56801 57335 56853
rect 57279 56799 57335 56801
rect 27788 55053 27844 55055
rect 27788 55001 27790 55053
rect 27790 55001 27842 55053
rect 27842 55001 27844 55053
rect 27788 54999 27844 55001
rect 27999 55053 28055 55055
rect 27999 55001 28001 55053
rect 28001 55001 28053 55053
rect 28053 55001 28055 55053
rect 27999 54999 28055 55001
rect 28210 55053 28266 55055
rect 28210 55001 28212 55053
rect 28212 55001 28264 55053
rect 28264 55001 28266 55053
rect 28210 54999 28266 55001
rect 28421 55053 28477 55055
rect 28421 55001 28423 55053
rect 28423 55001 28475 55053
rect 28475 55001 28477 55053
rect 28421 54999 28477 55001
rect 28632 55053 28688 55055
rect 28632 55001 28634 55053
rect 28634 55001 28686 55053
rect 28686 55001 28688 55053
rect 28632 54999 28688 55001
rect 28843 55053 28899 55055
rect 28843 55001 28845 55053
rect 28845 55001 28897 55053
rect 28897 55001 28899 55053
rect 28843 54999 28899 55001
rect 29054 55053 29110 55055
rect 29054 55001 29056 55053
rect 29056 55001 29108 55053
rect 29108 55001 29110 55053
rect 29054 54999 29110 55001
rect 56013 55053 56069 55055
rect 56013 55001 56015 55053
rect 56015 55001 56067 55053
rect 56067 55001 56069 55053
rect 56013 54999 56069 55001
rect 56224 55053 56280 55055
rect 56224 55001 56226 55053
rect 56226 55001 56278 55053
rect 56278 55001 56280 55053
rect 56224 54999 56280 55001
rect 56435 55053 56491 55055
rect 56435 55001 56437 55053
rect 56437 55001 56489 55053
rect 56489 55001 56491 55053
rect 56435 54999 56491 55001
rect 56646 55053 56702 55055
rect 56646 55001 56648 55053
rect 56648 55001 56700 55053
rect 56700 55001 56702 55053
rect 56646 54999 56702 55001
rect 56857 55053 56913 55055
rect 56857 55001 56859 55053
rect 56859 55001 56911 55053
rect 56911 55001 56913 55053
rect 56857 54999 56913 55001
rect 57068 55053 57124 55055
rect 57068 55001 57070 55053
rect 57070 55001 57122 55053
rect 57122 55001 57124 55053
rect 57068 54999 57124 55001
rect 57279 55053 57335 55055
rect 57279 55001 57281 55053
rect 57281 55001 57333 55053
rect 57333 55001 57335 55053
rect 57279 54999 57335 55001
rect 27788 53253 27844 53255
rect 27788 53201 27790 53253
rect 27790 53201 27842 53253
rect 27842 53201 27844 53253
rect 27788 53199 27844 53201
rect 27999 53253 28055 53255
rect 27999 53201 28001 53253
rect 28001 53201 28053 53253
rect 28053 53201 28055 53253
rect 27999 53199 28055 53201
rect 28210 53253 28266 53255
rect 28210 53201 28212 53253
rect 28212 53201 28264 53253
rect 28264 53201 28266 53253
rect 28210 53199 28266 53201
rect 28421 53253 28477 53255
rect 28421 53201 28423 53253
rect 28423 53201 28475 53253
rect 28475 53201 28477 53253
rect 28421 53199 28477 53201
rect 28632 53253 28688 53255
rect 28632 53201 28634 53253
rect 28634 53201 28686 53253
rect 28686 53201 28688 53253
rect 28632 53199 28688 53201
rect 28843 53253 28899 53255
rect 28843 53201 28845 53253
rect 28845 53201 28897 53253
rect 28897 53201 28899 53253
rect 28843 53199 28899 53201
rect 29054 53253 29110 53255
rect 29054 53201 29056 53253
rect 29056 53201 29108 53253
rect 29108 53201 29110 53253
rect 29054 53199 29110 53201
rect 56013 53253 56069 53255
rect 56013 53201 56015 53253
rect 56015 53201 56067 53253
rect 56067 53201 56069 53253
rect 56013 53199 56069 53201
rect 56224 53253 56280 53255
rect 56224 53201 56226 53253
rect 56226 53201 56278 53253
rect 56278 53201 56280 53253
rect 56224 53199 56280 53201
rect 56435 53253 56491 53255
rect 56435 53201 56437 53253
rect 56437 53201 56489 53253
rect 56489 53201 56491 53253
rect 56435 53199 56491 53201
rect 56646 53253 56702 53255
rect 56646 53201 56648 53253
rect 56648 53201 56700 53253
rect 56700 53201 56702 53253
rect 56646 53199 56702 53201
rect 56857 53253 56913 53255
rect 56857 53201 56859 53253
rect 56859 53201 56911 53253
rect 56911 53201 56913 53253
rect 56857 53199 56913 53201
rect 57068 53253 57124 53255
rect 57068 53201 57070 53253
rect 57070 53201 57122 53253
rect 57122 53201 57124 53253
rect 57068 53199 57124 53201
rect 57279 53253 57335 53255
rect 57279 53201 57281 53253
rect 57281 53201 57333 53253
rect 57333 53201 57335 53253
rect 57279 53199 57335 53201
rect 27788 51453 27844 51455
rect 27788 51401 27790 51453
rect 27790 51401 27842 51453
rect 27842 51401 27844 51453
rect 27788 51399 27844 51401
rect 27999 51453 28055 51455
rect 27999 51401 28001 51453
rect 28001 51401 28053 51453
rect 28053 51401 28055 51453
rect 27999 51399 28055 51401
rect 28210 51453 28266 51455
rect 28210 51401 28212 51453
rect 28212 51401 28264 51453
rect 28264 51401 28266 51453
rect 28210 51399 28266 51401
rect 28421 51453 28477 51455
rect 28421 51401 28423 51453
rect 28423 51401 28475 51453
rect 28475 51401 28477 51453
rect 28421 51399 28477 51401
rect 28632 51453 28688 51455
rect 28632 51401 28634 51453
rect 28634 51401 28686 51453
rect 28686 51401 28688 51453
rect 28632 51399 28688 51401
rect 28843 51453 28899 51455
rect 28843 51401 28845 51453
rect 28845 51401 28897 51453
rect 28897 51401 28899 51453
rect 28843 51399 28899 51401
rect 29054 51453 29110 51455
rect 29054 51401 29056 51453
rect 29056 51401 29108 51453
rect 29108 51401 29110 51453
rect 29054 51399 29110 51401
rect 56013 51453 56069 51455
rect 56013 51401 56015 51453
rect 56015 51401 56067 51453
rect 56067 51401 56069 51453
rect 56013 51399 56069 51401
rect 56224 51453 56280 51455
rect 56224 51401 56226 51453
rect 56226 51401 56278 51453
rect 56278 51401 56280 51453
rect 56224 51399 56280 51401
rect 56435 51453 56491 51455
rect 56435 51401 56437 51453
rect 56437 51401 56489 51453
rect 56489 51401 56491 51453
rect 56435 51399 56491 51401
rect 56646 51453 56702 51455
rect 56646 51401 56648 51453
rect 56648 51401 56700 51453
rect 56700 51401 56702 51453
rect 56646 51399 56702 51401
rect 56857 51453 56913 51455
rect 56857 51401 56859 51453
rect 56859 51401 56911 51453
rect 56911 51401 56913 51453
rect 56857 51399 56913 51401
rect 57068 51453 57124 51455
rect 57068 51401 57070 51453
rect 57070 51401 57122 51453
rect 57122 51401 57124 51453
rect 57068 51399 57124 51401
rect 57279 51453 57335 51455
rect 57279 51401 57281 51453
rect 57281 51401 57333 51453
rect 57333 51401 57335 51453
rect 57279 51399 57335 51401
rect 27788 49653 27844 49655
rect 27788 49601 27790 49653
rect 27790 49601 27842 49653
rect 27842 49601 27844 49653
rect 27788 49599 27844 49601
rect 27999 49653 28055 49655
rect 27999 49601 28001 49653
rect 28001 49601 28053 49653
rect 28053 49601 28055 49653
rect 27999 49599 28055 49601
rect 28210 49653 28266 49655
rect 28210 49601 28212 49653
rect 28212 49601 28264 49653
rect 28264 49601 28266 49653
rect 28210 49599 28266 49601
rect 28421 49653 28477 49655
rect 28421 49601 28423 49653
rect 28423 49601 28475 49653
rect 28475 49601 28477 49653
rect 28421 49599 28477 49601
rect 28632 49653 28688 49655
rect 28632 49601 28634 49653
rect 28634 49601 28686 49653
rect 28686 49601 28688 49653
rect 28632 49599 28688 49601
rect 28843 49653 28899 49655
rect 28843 49601 28845 49653
rect 28845 49601 28897 49653
rect 28897 49601 28899 49653
rect 28843 49599 28899 49601
rect 29054 49653 29110 49655
rect 29054 49601 29056 49653
rect 29056 49601 29108 49653
rect 29108 49601 29110 49653
rect 29054 49599 29110 49601
rect 56013 49653 56069 49655
rect 56013 49601 56015 49653
rect 56015 49601 56067 49653
rect 56067 49601 56069 49653
rect 56013 49599 56069 49601
rect 56224 49653 56280 49655
rect 56224 49601 56226 49653
rect 56226 49601 56278 49653
rect 56278 49601 56280 49653
rect 56224 49599 56280 49601
rect 56435 49653 56491 49655
rect 56435 49601 56437 49653
rect 56437 49601 56489 49653
rect 56489 49601 56491 49653
rect 56435 49599 56491 49601
rect 56646 49653 56702 49655
rect 56646 49601 56648 49653
rect 56648 49601 56700 49653
rect 56700 49601 56702 49653
rect 56646 49599 56702 49601
rect 56857 49653 56913 49655
rect 56857 49601 56859 49653
rect 56859 49601 56911 49653
rect 56911 49601 56913 49653
rect 56857 49599 56913 49601
rect 57068 49653 57124 49655
rect 57068 49601 57070 49653
rect 57070 49601 57122 49653
rect 57122 49601 57124 49653
rect 57068 49599 57124 49601
rect 57279 49653 57335 49655
rect 57279 49601 57281 49653
rect 57281 49601 57333 49653
rect 57333 49601 57335 49653
rect 57279 49599 57335 49601
rect 27788 47853 27844 47855
rect 27788 47801 27790 47853
rect 27790 47801 27842 47853
rect 27842 47801 27844 47853
rect 27788 47799 27844 47801
rect 27999 47853 28055 47855
rect 27999 47801 28001 47853
rect 28001 47801 28053 47853
rect 28053 47801 28055 47853
rect 27999 47799 28055 47801
rect 28210 47853 28266 47855
rect 28210 47801 28212 47853
rect 28212 47801 28264 47853
rect 28264 47801 28266 47853
rect 28210 47799 28266 47801
rect 28421 47853 28477 47855
rect 28421 47801 28423 47853
rect 28423 47801 28475 47853
rect 28475 47801 28477 47853
rect 28421 47799 28477 47801
rect 28632 47853 28688 47855
rect 28632 47801 28634 47853
rect 28634 47801 28686 47853
rect 28686 47801 28688 47853
rect 28632 47799 28688 47801
rect 28843 47853 28899 47855
rect 28843 47801 28845 47853
rect 28845 47801 28897 47853
rect 28897 47801 28899 47853
rect 28843 47799 28899 47801
rect 29054 47853 29110 47855
rect 29054 47801 29056 47853
rect 29056 47801 29108 47853
rect 29108 47801 29110 47853
rect 29054 47799 29110 47801
rect 56013 47853 56069 47855
rect 56013 47801 56015 47853
rect 56015 47801 56067 47853
rect 56067 47801 56069 47853
rect 56013 47799 56069 47801
rect 56224 47853 56280 47855
rect 56224 47801 56226 47853
rect 56226 47801 56278 47853
rect 56278 47801 56280 47853
rect 56224 47799 56280 47801
rect 56435 47853 56491 47855
rect 56435 47801 56437 47853
rect 56437 47801 56489 47853
rect 56489 47801 56491 47853
rect 56435 47799 56491 47801
rect 56646 47853 56702 47855
rect 56646 47801 56648 47853
rect 56648 47801 56700 47853
rect 56700 47801 56702 47853
rect 56646 47799 56702 47801
rect 56857 47853 56913 47855
rect 56857 47801 56859 47853
rect 56859 47801 56911 47853
rect 56911 47801 56913 47853
rect 56857 47799 56913 47801
rect 57068 47853 57124 47855
rect 57068 47801 57070 47853
rect 57070 47801 57122 47853
rect 57122 47801 57124 47853
rect 57068 47799 57124 47801
rect 57279 47853 57335 47855
rect 57279 47801 57281 47853
rect 57281 47801 57333 47853
rect 57333 47801 57335 47853
rect 57279 47799 57335 47801
rect 27788 46053 27844 46055
rect 27788 46001 27790 46053
rect 27790 46001 27842 46053
rect 27842 46001 27844 46053
rect 27788 45999 27844 46001
rect 27999 46053 28055 46055
rect 27999 46001 28001 46053
rect 28001 46001 28053 46053
rect 28053 46001 28055 46053
rect 27999 45999 28055 46001
rect 28210 46053 28266 46055
rect 28210 46001 28212 46053
rect 28212 46001 28264 46053
rect 28264 46001 28266 46053
rect 28210 45999 28266 46001
rect 28421 46053 28477 46055
rect 28421 46001 28423 46053
rect 28423 46001 28475 46053
rect 28475 46001 28477 46053
rect 28421 45999 28477 46001
rect 28632 46053 28688 46055
rect 28632 46001 28634 46053
rect 28634 46001 28686 46053
rect 28686 46001 28688 46053
rect 28632 45999 28688 46001
rect 28843 46053 28899 46055
rect 28843 46001 28845 46053
rect 28845 46001 28897 46053
rect 28897 46001 28899 46053
rect 28843 45999 28899 46001
rect 29054 46053 29110 46055
rect 29054 46001 29056 46053
rect 29056 46001 29108 46053
rect 29108 46001 29110 46053
rect 29054 45999 29110 46001
rect 56013 46053 56069 46055
rect 56013 46001 56015 46053
rect 56015 46001 56067 46053
rect 56067 46001 56069 46053
rect 56013 45999 56069 46001
rect 56224 46053 56280 46055
rect 56224 46001 56226 46053
rect 56226 46001 56278 46053
rect 56278 46001 56280 46053
rect 56224 45999 56280 46001
rect 56435 46053 56491 46055
rect 56435 46001 56437 46053
rect 56437 46001 56489 46053
rect 56489 46001 56491 46053
rect 56435 45999 56491 46001
rect 56646 46053 56702 46055
rect 56646 46001 56648 46053
rect 56648 46001 56700 46053
rect 56700 46001 56702 46053
rect 56646 45999 56702 46001
rect 56857 46053 56913 46055
rect 56857 46001 56859 46053
rect 56859 46001 56911 46053
rect 56911 46001 56913 46053
rect 56857 45999 56913 46001
rect 57068 46053 57124 46055
rect 57068 46001 57070 46053
rect 57070 46001 57122 46053
rect 57122 46001 57124 46053
rect 57068 45999 57124 46001
rect 57279 46053 57335 46055
rect 57279 46001 57281 46053
rect 57281 46001 57333 46053
rect 57333 46001 57335 46053
rect 57279 45999 57335 46001
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 26859 32032 26915 32088
rect 27071 32032 27127 32088
rect 26859 31814 26915 31870
rect 27071 31814 27127 31870
rect 26859 31596 26915 31652
rect 27071 31596 27127 31652
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 26924 20410 27084 20570
rect 26924 20066 27084 20226
rect 26465 19532 26625 19692
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 51766 9811 51822 9971
rect 49897 8897 50057 8953
rect 27474 7479 27530 7535
rect 27686 7479 27742 7535
rect 27474 7261 27530 7317
rect 27686 7261 27742 7317
rect 27474 7043 27530 7099
rect 27686 7043 27742 7099
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 5483 26915 5539
rect 27071 5483 27127 5539
rect 26859 5265 26915 5321
rect 27071 5265 27127 5321
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 43800 2994 43960 3050
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 32032 58052 32088
rect 58208 32032 58264 32088
rect 57996 31814 58052 31870
rect 58208 31814 58264 31870
rect 57996 31596 58052 31652
rect 58208 31596 58264 31652
rect 58048 20410 58208 20570
rect 58048 20066 58208 20226
rect 57996 5483 58052 5539
rect 58208 5483 58264 5539
rect 57996 5265 58052 5321
rect 58208 5265 58264 5321
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
<< metal3 >>
rect 1401 96176 2401 96976
rect 2626 96368 3626 96976
rect 4137 96176 5137 96976
rect 5362 96368 6362 96976
rect 6801 96176 7801 96976
rect 8026 96368 9026 96976
rect 9537 96176 10537 96976
rect 10762 96368 11762 96976
rect 12201 96176 13201 96976
rect 13426 96368 14426 96976
rect 14937 96176 15937 96976
rect 16162 96368 17162 96976
rect 17601 96176 18601 96976
rect 18826 96368 19826 96976
rect 20653 96176 21653 96976
rect 22258 96368 23258 96976
rect 23483 96176 24483 96976
rect 25158 96368 26158 96976
rect 26572 96176 27572 96976
rect 27877 96368 28877 96976
rect 29273 96368 30273 96976
rect 30710 96176 31710 96976
rect 32381 96368 33381 96976
rect 34024 96368 35024 96976
rect 35415 96176 36415 96976
rect 36948 96368 37948 96976
rect 38585 96176 39585 96976
rect 39882 96368 40882 96976
rect 41230 96176 42230 96976
rect 42430 96368 43430 96976
rect 43713 96368 44713 96976
rect 45069 96176 46069 96976
rect 46313 96176 47313 96976
rect 47538 96368 48538 96976
rect 48901 96176 49901 96976
rect 50465 96368 51465 96976
rect 52569 96176 53569 96976
rect 54262 96176 55262 96976
rect 55990 96368 56990 96976
rect 57547 96176 58547 96976
rect 58791 96368 59791 96976
rect 60977 96176 61977 96976
rect 62202 96368 63202 96976
rect 63713 96176 64713 96976
rect 64938 96368 65938 96976
rect 66377 96176 67377 96976
rect 67602 96368 68602 96976
rect 69113 96176 70113 96976
rect 70338 96368 71338 96976
rect 71777 96176 72777 96976
rect 73002 96368 74002 96976
rect 74513 96176 75513 96976
rect 75738 96368 76738 96976
rect 77177 96176 78177 96976
rect 78402 96368 79402 96976
rect 80229 96176 81229 96976
rect 81834 96368 82834 96976
rect 83059 96176 84059 96976
rect 84666 96176 85666 96976
rect 0 95176 86372 96176
rect 0 94776 1014 94976
rect 25376 94776 25948 94785
rect 58855 94776 59427 94785
rect 85358 94776 86372 94976
rect 0 94728 27272 94776
rect 58855 94728 86372 94776
rect 0 94655 86372 94728
rect 0 94599 27788 94655
rect 27844 94599 27999 94655
rect 28055 94599 28210 94655
rect 28266 94599 28421 94655
rect 28477 94599 28632 94655
rect 28688 94599 28843 94655
rect 28899 94599 29054 94655
rect 29110 94599 56013 94655
rect 56069 94599 56224 94655
rect 56280 94599 56435 94655
rect 56491 94599 56646 94655
rect 56702 94599 56857 94655
rect 56913 94599 57068 94655
rect 57124 94599 57279 94655
rect 57335 94599 86372 94655
rect 0 94527 86372 94599
rect 0 94476 27272 94527
rect 30402 94526 54622 94527
rect 58855 94476 86372 94527
rect 0 94276 1014 94476
rect 25376 94461 25948 94476
rect 58855 94461 59427 94476
rect 85358 94276 86372 94476
rect 0 93376 1706 94076
rect 56271 94066 61644 94268
rect 84666 93376 86372 94076
rect 0 92976 1014 93176
rect 85358 92976 86372 93176
rect 0 92928 27272 92976
rect 59421 92928 86372 92976
rect 0 92855 86372 92928
rect 0 92799 27788 92855
rect 27844 92799 27999 92855
rect 28055 92799 28210 92855
rect 28266 92799 28421 92855
rect 28477 92799 28632 92855
rect 28688 92799 28843 92855
rect 28899 92799 29054 92855
rect 29110 92799 56013 92855
rect 56069 92799 56224 92855
rect 56280 92799 56435 92855
rect 56491 92799 56646 92855
rect 56702 92799 56857 92855
rect 56913 92799 57068 92855
rect 57124 92799 57279 92855
rect 57335 92799 86372 92855
rect 0 92727 86372 92799
rect 0 92676 27272 92727
rect 30403 92726 54622 92727
rect 59421 92676 86372 92727
rect 0 92476 1014 92676
rect 85358 92476 86372 92676
rect 0 91576 1706 92276
rect 84666 91576 86372 92276
rect 0 91176 1014 91376
rect 85358 91176 86372 91376
rect 0 91128 27272 91176
rect 59421 91128 86372 91176
rect 0 91055 86372 91128
rect 0 90999 27788 91055
rect 27844 90999 27999 91055
rect 28055 90999 28210 91055
rect 28266 90999 28421 91055
rect 28477 90999 28632 91055
rect 28688 90999 28843 91055
rect 28899 90999 29054 91055
rect 29110 90999 56013 91055
rect 56069 90999 56224 91055
rect 56280 90999 56435 91055
rect 56491 90999 56646 91055
rect 56702 90999 56857 91055
rect 56913 90999 57068 91055
rect 57124 90999 57279 91055
rect 57335 90999 86372 91055
rect 0 90927 86372 90999
rect 0 90876 27272 90927
rect 30403 90926 54622 90927
rect 59421 90876 86372 90927
rect 0 90676 1014 90876
rect 85358 90676 86372 90876
rect 0 89776 1706 90476
rect 84666 89776 86372 90476
rect 0 89376 1014 89576
rect 85358 89376 86372 89576
rect 0 89328 27272 89376
rect 59421 89328 86372 89376
rect 0 89255 86372 89328
rect 0 89199 27788 89255
rect 27844 89199 27999 89255
rect 28055 89199 28210 89255
rect 28266 89199 28421 89255
rect 28477 89199 28632 89255
rect 28688 89199 28843 89255
rect 28899 89199 29054 89255
rect 29110 89199 56013 89255
rect 56069 89199 56224 89255
rect 56280 89199 56435 89255
rect 56491 89199 56646 89255
rect 56702 89199 56857 89255
rect 56913 89199 57068 89255
rect 57124 89199 57279 89255
rect 57335 89199 86372 89255
rect 0 89127 86372 89199
rect 0 89076 27272 89127
rect 30403 89126 54622 89127
rect 59421 89076 86372 89127
rect 0 88876 1014 89076
rect 85358 88876 86372 89076
rect 0 87976 1706 88676
rect 84666 87976 86372 88676
rect 0 87576 1014 87776
rect 85358 87576 86372 87776
rect 0 87528 27272 87576
rect 59421 87528 86372 87576
rect 0 87455 86372 87528
rect 0 87399 27788 87455
rect 27844 87399 27999 87455
rect 28055 87399 28210 87455
rect 28266 87399 28421 87455
rect 28477 87399 28632 87455
rect 28688 87399 28843 87455
rect 28899 87399 29054 87455
rect 29110 87399 56013 87455
rect 56069 87399 56224 87455
rect 56280 87399 56435 87455
rect 56491 87399 56646 87455
rect 56702 87399 56857 87455
rect 56913 87399 57068 87455
rect 57124 87399 57279 87455
rect 57335 87399 86372 87455
rect 0 87327 86372 87399
rect 0 87276 27272 87327
rect 30403 87326 54622 87327
rect 59421 87276 86372 87327
rect 0 87076 1014 87276
rect 85358 87076 86372 87276
rect 0 86176 1706 86876
rect 84666 86176 86372 86876
rect 0 85776 1014 85976
rect 85358 85776 86372 85976
rect 0 85728 27272 85776
rect 59421 85728 86372 85776
rect 0 85655 86372 85728
rect 0 85599 27788 85655
rect 27844 85599 27999 85655
rect 28055 85599 28210 85655
rect 28266 85599 28421 85655
rect 28477 85599 28632 85655
rect 28688 85599 28843 85655
rect 28899 85599 29054 85655
rect 29110 85599 56013 85655
rect 56069 85599 56224 85655
rect 56280 85599 56435 85655
rect 56491 85599 56646 85655
rect 56702 85599 56857 85655
rect 56913 85599 57068 85655
rect 57124 85599 57279 85655
rect 57335 85599 86372 85655
rect 0 85527 86372 85599
rect 0 85476 27272 85527
rect 30403 85526 54622 85527
rect 59421 85476 86372 85527
rect 0 85276 1014 85476
rect 85358 85276 86372 85476
rect 0 84376 1706 85076
rect 84666 84376 86372 85076
rect 0 83976 1014 84176
rect 85358 83976 86372 84176
rect 0 83928 27272 83976
rect 59421 83928 86372 83976
rect 0 83855 86372 83928
rect 0 83799 27788 83855
rect 27844 83799 27999 83855
rect 28055 83799 28210 83855
rect 28266 83799 28421 83855
rect 28477 83799 28632 83855
rect 28688 83799 28843 83855
rect 28899 83799 29054 83855
rect 29110 83799 56013 83855
rect 56069 83799 56224 83855
rect 56280 83799 56435 83855
rect 56491 83799 56646 83855
rect 56702 83799 56857 83855
rect 56913 83799 57068 83855
rect 57124 83799 57279 83855
rect 57335 83799 86372 83855
rect 0 83727 86372 83799
rect 0 83676 27272 83727
rect 30403 83726 54622 83727
rect 59421 83676 86372 83727
rect 0 83476 1014 83676
rect 85358 83476 86372 83676
rect 0 82576 1706 83276
rect 84666 82576 86372 83276
rect 0 82176 1014 82376
rect 85358 82176 86372 82376
rect 0 82128 27272 82176
rect 59421 82128 86372 82176
rect 0 82055 86372 82128
rect 0 81999 27788 82055
rect 27844 81999 27999 82055
rect 28055 81999 28210 82055
rect 28266 81999 28421 82055
rect 28477 81999 28632 82055
rect 28688 81999 28843 82055
rect 28899 81999 29054 82055
rect 29110 81999 56013 82055
rect 56069 81999 56224 82055
rect 56280 81999 56435 82055
rect 56491 81999 56646 82055
rect 56702 81999 56857 82055
rect 56913 81999 57068 82055
rect 57124 81999 57279 82055
rect 57335 81999 86372 82055
rect 0 81927 86372 81999
rect 0 81876 27272 81927
rect 30403 81926 54622 81927
rect 59421 81876 86372 81927
rect 0 81676 1014 81876
rect 85358 81676 86372 81876
rect 0 80776 1706 81476
rect 84666 80776 86372 81476
rect 0 80376 1014 80576
rect 85358 80376 86372 80576
rect 0 80328 27272 80376
rect 59421 80328 86372 80376
rect 0 80255 86372 80328
rect 0 80199 27788 80255
rect 27844 80199 27999 80255
rect 28055 80199 28210 80255
rect 28266 80199 28421 80255
rect 28477 80199 28632 80255
rect 28688 80199 28843 80255
rect 28899 80199 29054 80255
rect 29110 80199 56013 80255
rect 56069 80199 56224 80255
rect 56280 80199 56435 80255
rect 56491 80199 56646 80255
rect 56702 80199 56857 80255
rect 56913 80199 57068 80255
rect 57124 80199 57279 80255
rect 57335 80199 86372 80255
rect 0 80127 86372 80199
rect 0 80076 27272 80127
rect 30403 80126 54622 80127
rect 59421 80076 86372 80127
rect 0 79876 1014 80076
rect 85358 79876 86372 80076
rect 0 78976 1706 79676
rect 84666 78976 86372 79676
rect 0 78576 1014 78776
rect 85358 78576 86372 78776
rect 0 78528 27272 78576
rect 59421 78528 86372 78576
rect 0 78455 86372 78528
rect 0 78399 27788 78455
rect 27844 78399 27999 78455
rect 28055 78399 28210 78455
rect 28266 78399 28421 78455
rect 28477 78399 28632 78455
rect 28688 78399 28843 78455
rect 28899 78399 29054 78455
rect 29110 78399 56013 78455
rect 56069 78399 56224 78455
rect 56280 78399 56435 78455
rect 56491 78399 56646 78455
rect 56702 78399 56857 78455
rect 56913 78399 57068 78455
rect 57124 78399 57279 78455
rect 57335 78399 86372 78455
rect 0 78327 86372 78399
rect 0 78276 27272 78327
rect 30403 78326 54622 78327
rect 59421 78276 86372 78327
rect 0 78076 1014 78276
rect 85358 78076 86372 78276
rect 0 77176 1706 77876
rect 84666 77176 86372 77876
rect 0 76776 1014 76976
rect 85358 76776 86372 76976
rect 0 76728 27272 76776
rect 59421 76728 86372 76776
rect 0 76655 86372 76728
rect 0 76599 27788 76655
rect 27844 76599 27999 76655
rect 28055 76599 28210 76655
rect 28266 76599 28421 76655
rect 28477 76599 28632 76655
rect 28688 76599 28843 76655
rect 28899 76599 29054 76655
rect 29110 76599 56013 76655
rect 56069 76599 56224 76655
rect 56280 76599 56435 76655
rect 56491 76599 56646 76655
rect 56702 76599 56857 76655
rect 56913 76599 57068 76655
rect 57124 76599 57279 76655
rect 57335 76599 86372 76655
rect 0 76527 86372 76599
rect 0 76476 27272 76527
rect 30403 76526 54622 76527
rect 59421 76476 86372 76527
rect 0 76276 1014 76476
rect 85358 76276 86372 76476
rect 0 75376 1706 76076
rect 84666 75376 86372 76076
rect 0 74976 1014 75176
rect 85358 74976 86372 75176
rect 0 74928 27272 74976
rect 59421 74928 86372 74976
rect 0 74855 86372 74928
rect 0 74799 27788 74855
rect 27844 74799 27999 74855
rect 28055 74799 28210 74855
rect 28266 74799 28421 74855
rect 28477 74799 28632 74855
rect 28688 74799 28843 74855
rect 28899 74799 29054 74855
rect 29110 74799 56013 74855
rect 56069 74799 56224 74855
rect 56280 74799 56435 74855
rect 56491 74799 56646 74855
rect 56702 74799 56857 74855
rect 56913 74799 57068 74855
rect 57124 74799 57279 74855
rect 57335 74799 86372 74855
rect 0 74727 86372 74799
rect 0 74676 27272 74727
rect 30403 74726 54622 74727
rect 59421 74676 86372 74727
rect 0 74476 1014 74676
rect 85358 74476 86372 74676
rect 0 73576 1706 74276
rect 84666 73576 86372 74276
rect 0 73176 1014 73376
rect 85358 73176 86372 73376
rect 0 73128 27272 73176
rect 59421 73128 86372 73176
rect 0 73055 86372 73128
rect 0 72999 27788 73055
rect 27844 72999 27999 73055
rect 28055 72999 28210 73055
rect 28266 72999 28421 73055
rect 28477 72999 28632 73055
rect 28688 72999 28843 73055
rect 28899 72999 29054 73055
rect 29110 72999 56013 73055
rect 56069 72999 56224 73055
rect 56280 72999 56435 73055
rect 56491 72999 56646 73055
rect 56702 72999 56857 73055
rect 56913 72999 57068 73055
rect 57124 72999 57279 73055
rect 57335 72999 86372 73055
rect 0 72927 86372 72999
rect 0 72876 27272 72927
rect 30403 72926 54622 72927
rect 59421 72876 86372 72927
rect 0 72676 1014 72876
rect 85358 72676 86372 72876
rect 0 71776 1706 72476
rect 84666 71776 86372 72476
rect 0 71376 1014 71576
rect 85358 71376 86372 71576
rect 0 71328 27272 71376
rect 59421 71328 86372 71376
rect 0 71255 86372 71328
rect 0 71199 27788 71255
rect 27844 71199 27999 71255
rect 28055 71199 28210 71255
rect 28266 71199 28421 71255
rect 28477 71199 28632 71255
rect 28688 71199 28843 71255
rect 28899 71199 29054 71255
rect 29110 71199 56013 71255
rect 56069 71199 56224 71255
rect 56280 71199 56435 71255
rect 56491 71199 56646 71255
rect 56702 71199 56857 71255
rect 56913 71199 57068 71255
rect 57124 71199 57279 71255
rect 57335 71199 86372 71255
rect 0 71127 86372 71199
rect 0 71076 27272 71127
rect 30403 71126 54622 71127
rect 59421 71076 86372 71127
rect 0 70876 1014 71076
rect 85358 70876 86372 71076
rect 0 69976 1706 70676
rect 84666 69976 86372 70676
rect 0 69576 1014 69776
rect 85358 69576 86372 69776
rect 0 69528 27272 69576
rect 59421 69528 86372 69576
rect 0 69455 86372 69528
rect 0 69399 27788 69455
rect 27844 69399 27999 69455
rect 28055 69399 28210 69455
rect 28266 69399 28421 69455
rect 28477 69399 28632 69455
rect 28688 69399 28843 69455
rect 28899 69399 29054 69455
rect 29110 69399 56013 69455
rect 56069 69399 56224 69455
rect 56280 69399 56435 69455
rect 56491 69399 56646 69455
rect 56702 69399 56857 69455
rect 56913 69399 57068 69455
rect 57124 69399 57279 69455
rect 57335 69399 86372 69455
rect 0 69327 86372 69399
rect 0 69276 27272 69327
rect 30403 69326 54622 69327
rect 59421 69276 86372 69327
rect 0 69076 1014 69276
rect 85358 69076 86372 69276
rect 0 68176 1706 68876
rect 84666 68176 86372 68876
rect 0 67776 1014 67976
rect 85358 67776 86372 67976
rect 0 67728 27272 67776
rect 59421 67728 86372 67776
rect 0 67655 86372 67728
rect 0 67599 27788 67655
rect 27844 67599 27999 67655
rect 28055 67599 28210 67655
rect 28266 67599 28421 67655
rect 28477 67599 28632 67655
rect 28688 67599 28843 67655
rect 28899 67599 29054 67655
rect 29110 67599 56013 67655
rect 56069 67599 56224 67655
rect 56280 67599 56435 67655
rect 56491 67599 56646 67655
rect 56702 67599 56857 67655
rect 56913 67599 57068 67655
rect 57124 67599 57279 67655
rect 57335 67599 86372 67655
rect 0 67527 86372 67599
rect 0 67476 27272 67527
rect 30403 67526 54622 67527
rect 59421 67476 86372 67527
rect 0 67276 1014 67476
rect 85358 67276 86372 67476
rect 0 66376 1706 67076
rect 84666 66376 86372 67076
rect 0 65976 1014 66176
rect 85358 65976 86372 66176
rect 0 65928 27272 65976
rect 59421 65928 86372 65976
rect 0 65855 86372 65928
rect 0 65799 27788 65855
rect 27844 65799 27999 65855
rect 28055 65799 28210 65855
rect 28266 65799 28421 65855
rect 28477 65799 28632 65855
rect 28688 65799 28843 65855
rect 28899 65799 29054 65855
rect 29110 65799 56013 65855
rect 56069 65799 56224 65855
rect 56280 65799 56435 65855
rect 56491 65799 56646 65855
rect 56702 65799 56857 65855
rect 56913 65799 57068 65855
rect 57124 65799 57279 65855
rect 57335 65799 86372 65855
rect 0 65727 86372 65799
rect 0 65676 27272 65727
rect 30403 65726 54622 65727
rect 59421 65676 86372 65727
rect 0 65476 1014 65676
rect 85358 65476 86372 65676
rect 0 64576 1706 65276
rect 84666 64576 86372 65276
rect 0 64176 1014 64376
rect 85358 64176 86372 64376
rect 0 64128 27272 64176
rect 59421 64128 86372 64176
rect 0 64055 86372 64128
rect 0 63999 27788 64055
rect 27844 63999 27999 64055
rect 28055 63999 28210 64055
rect 28266 63999 28421 64055
rect 28477 63999 28632 64055
rect 28688 63999 28843 64055
rect 28899 63999 29054 64055
rect 29110 63999 56013 64055
rect 56069 63999 56224 64055
rect 56280 63999 56435 64055
rect 56491 63999 56646 64055
rect 56702 63999 56857 64055
rect 56913 63999 57068 64055
rect 57124 63999 57279 64055
rect 57335 63999 86372 64055
rect 0 63927 86372 63999
rect 0 63876 27272 63927
rect 30403 63926 54622 63927
rect 59421 63876 86372 63927
rect 0 63676 1014 63876
rect 85358 63676 86372 63876
rect 0 62776 1706 63476
rect 84666 62776 86372 63476
rect 0 62376 1014 62576
rect 85358 62376 86372 62576
rect 0 62328 27272 62376
rect 59421 62328 86372 62376
rect 0 62255 86372 62328
rect 0 62199 27788 62255
rect 27844 62199 27999 62255
rect 28055 62199 28210 62255
rect 28266 62199 28421 62255
rect 28477 62199 28632 62255
rect 28688 62199 28843 62255
rect 28899 62199 29054 62255
rect 29110 62199 56013 62255
rect 56069 62199 56224 62255
rect 56280 62199 56435 62255
rect 56491 62199 56646 62255
rect 56702 62199 56857 62255
rect 56913 62199 57068 62255
rect 57124 62199 57279 62255
rect 57335 62199 86372 62255
rect 0 62127 86372 62199
rect 0 62076 27272 62127
rect 30403 62126 54622 62127
rect 59421 62076 86372 62127
rect 0 61876 1014 62076
rect 85358 61876 86372 62076
rect 0 60976 1706 61676
rect 84666 60976 86372 61676
rect 0 60576 1014 60776
rect 85358 60576 86372 60776
rect 0 60528 27272 60576
rect 59421 60528 86372 60576
rect 0 60455 86372 60528
rect 0 60399 27788 60455
rect 27844 60399 27999 60455
rect 28055 60399 28210 60455
rect 28266 60399 28421 60455
rect 28477 60399 28632 60455
rect 28688 60399 28843 60455
rect 28899 60399 29054 60455
rect 29110 60399 56013 60455
rect 56069 60399 56224 60455
rect 56280 60399 56435 60455
rect 56491 60399 56646 60455
rect 56702 60399 56857 60455
rect 56913 60399 57068 60455
rect 57124 60399 57279 60455
rect 57335 60399 86372 60455
rect 0 60327 86372 60399
rect 0 60276 27272 60327
rect 30403 60326 54622 60327
rect 59421 60276 86372 60327
rect 0 60076 1014 60276
rect 85358 60076 86372 60276
rect 0 59176 1706 59876
rect 84666 59176 86372 59876
rect 0 58776 1014 58976
rect 85358 58776 86372 58976
rect 0 58728 27272 58776
rect 59421 58728 86372 58776
rect 0 58655 86372 58728
rect 0 58599 27788 58655
rect 27844 58599 27999 58655
rect 28055 58599 28210 58655
rect 28266 58599 28421 58655
rect 28477 58599 28632 58655
rect 28688 58599 28843 58655
rect 28899 58599 29054 58655
rect 29110 58599 56013 58655
rect 56069 58599 56224 58655
rect 56280 58599 56435 58655
rect 56491 58599 56646 58655
rect 56702 58599 56857 58655
rect 56913 58599 57068 58655
rect 57124 58599 57279 58655
rect 57335 58599 86372 58655
rect 0 58527 86372 58599
rect 0 58476 27272 58527
rect 30403 58526 54622 58527
rect 59421 58476 86372 58527
rect 0 58276 1014 58476
rect 85358 58276 86372 58476
rect 0 57376 1706 58076
rect 84666 57376 86372 58076
rect 0 56976 1014 57176
rect 85358 56976 86372 57176
rect 0 56928 27272 56976
rect 59421 56928 86372 56976
rect 0 56855 86372 56928
rect 0 56799 27788 56855
rect 27844 56799 27999 56855
rect 28055 56799 28210 56855
rect 28266 56799 28421 56855
rect 28477 56799 28632 56855
rect 28688 56799 28843 56855
rect 28899 56799 29054 56855
rect 29110 56799 56013 56855
rect 56069 56799 56224 56855
rect 56280 56799 56435 56855
rect 56491 56799 56646 56855
rect 56702 56799 56857 56855
rect 56913 56799 57068 56855
rect 57124 56799 57279 56855
rect 57335 56799 86372 56855
rect 0 56727 86372 56799
rect 0 56676 27272 56727
rect 30403 56726 54622 56727
rect 59421 56676 86372 56727
rect 0 56476 1014 56676
rect 85358 56476 86372 56676
rect 0 55576 1706 56276
rect 84666 55576 86372 56276
rect 0 55176 1014 55376
rect 85358 55176 86372 55376
rect 0 55128 27272 55176
rect 59421 55128 86372 55176
rect 0 55055 86372 55128
rect 0 54999 27788 55055
rect 27844 54999 27999 55055
rect 28055 54999 28210 55055
rect 28266 54999 28421 55055
rect 28477 54999 28632 55055
rect 28688 54999 28843 55055
rect 28899 54999 29054 55055
rect 29110 54999 56013 55055
rect 56069 54999 56224 55055
rect 56280 54999 56435 55055
rect 56491 54999 56646 55055
rect 56702 54999 56857 55055
rect 56913 54999 57068 55055
rect 57124 54999 57279 55055
rect 57335 54999 86372 55055
rect 0 54927 86372 54999
rect 0 54876 27272 54927
rect 30403 54926 54622 54927
rect 59421 54876 86372 54927
rect 0 54676 1014 54876
rect 85358 54676 86372 54876
rect 0 53776 1706 54476
rect 84666 53776 86372 54476
rect 0 53376 1014 53576
rect 85358 53376 86372 53576
rect 0 53328 27272 53376
rect 59421 53328 86372 53376
rect 0 53255 86372 53328
rect 0 53199 27788 53255
rect 27844 53199 27999 53255
rect 28055 53199 28210 53255
rect 28266 53199 28421 53255
rect 28477 53199 28632 53255
rect 28688 53199 28843 53255
rect 28899 53199 29054 53255
rect 29110 53199 56013 53255
rect 56069 53199 56224 53255
rect 56280 53199 56435 53255
rect 56491 53199 56646 53255
rect 56702 53199 56857 53255
rect 56913 53199 57068 53255
rect 57124 53199 57279 53255
rect 57335 53199 86372 53255
rect 0 53127 86372 53199
rect 0 53076 27272 53127
rect 30403 53126 54622 53127
rect 59421 53076 86372 53127
rect 0 52876 1014 53076
rect 85358 52876 86372 53076
rect 0 51976 1706 52676
rect 84666 51976 86372 52676
rect 0 51576 1014 51776
rect 85358 51576 86372 51776
rect 0 51528 27272 51576
rect 59421 51528 86372 51576
rect 0 51455 86372 51528
rect 0 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 86372 51455
rect 0 51327 86372 51399
rect 0 51276 27272 51327
rect 30403 51326 54622 51327
rect 59421 51276 86372 51327
rect 0 51076 1014 51276
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49728 27272 49776
rect 59421 49728 86372 49776
rect 0 49655 86372 49728
rect 0 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 86372 49655
rect 0 49527 86372 49599
rect 0 49476 27272 49527
rect 30403 49526 54622 49527
rect 59421 49476 86372 49527
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47928 27272 47976
rect 59421 47928 86372 47976
rect 0 47855 86372 47928
rect 0 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 86372 47855
rect 0 47727 86372 47799
rect 0 47676 27272 47727
rect 30403 47726 54622 47727
rect 59421 47676 86372 47727
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46128 27272 46176
rect 59421 46128 86372 46176
rect 0 46055 86372 46128
rect 0 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 86372 46055
rect 0 45927 86372 45999
rect 0 45876 27272 45927
rect 30403 45926 54622 45927
rect 59421 45876 86372 45927
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44328 27272 44376
rect 59421 44328 86372 44376
rect 0 44255 86372 44328
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44127 86372 44199
rect 0 44076 27272 44127
rect 30403 44126 54622 44127
rect 59421 44076 86372 44127
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42528 27272 42576
rect 59421 42528 86372 42576
rect 0 42455 86372 42528
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42327 86372 42399
rect 0 42276 27272 42327
rect 30403 42326 54622 42327
rect 59421 42276 86372 42327
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40728 27272 40776
rect 59421 40728 86372 40776
rect 0 40655 86372 40728
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40527 86372 40599
rect 0 40476 27272 40527
rect 30403 40526 54622 40527
rect 59421 40476 86372 40527
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38928 27272 38976
rect 59421 38928 86372 38976
rect 0 38855 86372 38928
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38727 86372 38799
rect 0 38676 27272 38727
rect 30403 38726 54622 38727
rect 59421 38676 86372 38727
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37128 27272 37176
rect 59421 37128 86372 37176
rect 0 37055 86372 37128
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36927 86372 36999
rect 0 36876 27272 36927
rect 30403 36926 54622 36927
rect 59421 36876 86372 36927
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 35126 24917 35326
rect 0 35016 1014 35126
rect 0 34536 27830 35016
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 32318 27214 34124
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 83360 35298 86372 35326
rect 60460 35158 86372 35298
rect 83360 35126 86372 35158
rect 85358 35016 86372 35126
rect 58791 34536 86372 35016
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 33263
rect 56135 32311 57736 33263
rect 57908 32315 86372 34124
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 30443 28929 31352
rect 56186 30443 59524 31352
rect 26772 29714 58351 30105
rect 84666 29714 86372 32315
rect 0 29430 86372 29714
rect 0 28412 3011 28416
rect 0 26890 26070 28412
rect 26772 27382 58351 29430
rect 83361 28412 86372 28416
rect 58785 26890 86372 28412
rect 0 26799 27828 26890
rect 0 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 0 26581 27828 26743
rect 0 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 0 26435 27828 26525
rect 57295 26799 86372 26890
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 86372 26799
rect 57295 26581 86372 26743
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 86372 26581
rect 57295 26435 86372 26525
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 23425 26434 27828 26435
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23380 58348 24278
rect 84666 23380 86372 23938
rect 0 23370 86372 23380
rect 0 22938 27214 23370
rect 27387 22291 57681 23199
rect 57908 22938 86372 23370
rect 57908 22937 83763 22938
rect 27387 22282 27826 22291
rect 0 21827 27826 22282
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22282 57681 22291
rect 56078 21827 86372 22282
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61807 16784 86372 17730
rect 24111 16597 27828 16598
rect 0 15015 27828 16597
rect 46982 15015 86372 16784
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14936 51760 14966
rect 0 14491 47683 14936
rect 0 14329 45977 14491
rect 0 14328 24250 14329
rect 24047 14178 27214 14179
rect 0 13461 27214 14178
rect 0 12846 1706 13461
rect 24047 12934 27214 13461
rect 27387 13760 45977 14329
rect 57295 14328 86372 14968
rect 57295 14327 83763 14328
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13245 49775 13760
rect 29478 13243 49775 13245
rect 41493 13078 49775 13243
rect 50228 13461 86372 13866
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12570 34761 12846
rect 50228 12846 58421 13461
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12570 86372 12846
rect 0 12046 86372 12570
rect 0 12036 24250 12046
rect 26772 12036 86372 12046
rect 26772 12035 84999 12036
rect 26772 11844 58351 12035
rect 29478 11697 58351 11844
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 10176 27828 11491
rect 29478 10756 41516 11697
rect 61825 11491 86372 11493
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 23612 9942 29221 10030
rect 34741 9972 41516 10756
rect 42261 10740 86372 11491
rect 24047 9515 28729 9516
rect 0 9514 1014 9515
rect 2226 9514 28729 9515
rect 0 8154 28729 9514
rect 29133 9302 29221 9942
rect 41857 9502 51430 10420
rect 51750 10097 54952 10185
rect 57295 10176 86372 10740
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10030 54952 10097
rect 54864 9942 62145 10030
rect 51750 9801 51838 9811
rect 58688 9681 61743 9777
rect 57909 9515 62278 9516
rect 57909 9514 72434 9515
rect 72602 9514 83234 9515
rect 85358 9514 86372 9515
rect 29133 9214 41656 9302
rect 41568 8972 41656 9214
rect 41857 9165 55482 9502
rect 41568 8953 50067 8972
rect 41568 8897 49897 8953
rect 50057 8897 50067 8953
rect 41568 8884 50067 8897
rect 50922 8930 55482 9165
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6306 29058 6875
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 7596 57736 8930
rect 57909 8154 86372 9514
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7392 86372 7595
rect 34860 6984 86372 7392
rect 34860 6592 55482 6984
rect 61802 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6306 62747 6874
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5321 86372 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 86372 5321
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 61802 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60886 3420 86372 3524
rect 0 2854 1014 3420
rect 24169 3050 62588 3066
rect 24169 2994 43800 3050
rect 43960 2994 62588 3050
rect 24169 2978 62588 2994
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 512x8M8W_PWR_512x8m81  512x8M8W_PWR_512x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use GF018_512x8M8WM1_lef_512x8m81  GF018_512x8M8WM1_lef_512x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 0 0 86372 96976
use G_ring_512x8m81  G_ring_512x8m81_0
timestamp 1666464484
transform 1 0 282 0 1 0
box 0 0 85816 96702
use M1_PSUB4310591302010_512x8m81  M1_PSUB4310591302010_512x8m81_0
timestamp 1666464484
transform 1 0 53710 0 1 2781
box -2884 -1144 2884 1144
use M1_PSUB4310591302014_512x8m81  M1_PSUB4310591302014_512x8m81_0
timestamp 1666464484
transform 1 0 34404 0 1 2781
box -5784 -1144 5784 1144
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_0
timestamp 1666464484
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_1
timestamp 1666464484
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_2
timestamp 1666464484
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_3
timestamp 1666464484
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_4
timestamp 1666464484
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_5
timestamp 1666464484
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_6
timestamp 1666464484
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_7
timestamp 1666464484
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_8
timestamp 1666464484
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_9
timestamp 1666464484
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_10
timestamp 1666464484
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_11
timestamp 1666464484
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_12
timestamp 1666464484
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_13
timestamp 1666464484
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_14
timestamp 1666464484
transform 1 0 28449 0 1 92827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_15
timestamp 1666464484
transform 1 0 28449 0 1 91027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_16
timestamp 1666464484
transform 1 0 28449 0 1 89227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_17
timestamp 1666464484
transform 1 0 28449 0 1 87427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_18
timestamp 1666464484
transform 1 0 28449 0 1 85627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_19
timestamp 1666464484
transform 1 0 28449 0 1 83827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_20
timestamp 1666464484
transform 1 0 28449 0 1 82027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_21
timestamp 1666464484
transform 1 0 28449 0 1 80227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_22
timestamp 1666464484
transform 1 0 28449 0 1 78427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_23
timestamp 1666464484
transform 1 0 28449 0 1 76627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_24
timestamp 1666464484
transform 1 0 28449 0 1 74827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_25
timestamp 1666464484
transform 1 0 28449 0 1 73027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_26
timestamp 1666464484
transform 1 0 28449 0 1 71227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_27
timestamp 1666464484
transform 1 0 28449 0 1 69427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_28
timestamp 1666464484
transform 1 0 28449 0 1 67627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_29
timestamp 1666464484
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_30
timestamp 1666464484
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_31
timestamp 1666464484
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_32
timestamp 1666464484
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_33
timestamp 1666464484
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_34
timestamp 1666464484
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_35
timestamp 1666464484
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_36
timestamp 1666464484
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_37
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_38
timestamp 1666464484
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_39
timestamp 1666464484
transform 1 0 28449 0 1 94627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_40
timestamp 1666464484
transform 1 0 56674 0 1 87427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_41
timestamp 1666464484
transform 1 0 56674 0 1 89227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_42
timestamp 1666464484
transform 1 0 56674 0 1 91027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_43
timestamp 1666464484
transform 1 0 56674 0 1 92827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_44
timestamp 1666464484
transform 1 0 56674 0 1 94627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_45
timestamp 1666464484
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_46
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_47
timestamp 1666464484
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_48
timestamp 1666464484
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_49
timestamp 1666464484
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_50
timestamp 1666464484
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_51
timestamp 1666464484
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_52
timestamp 1666464484
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_53
timestamp 1666464484
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_54
timestamp 1666464484
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_55
timestamp 1666464484
transform 1 0 56674 0 1 67627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_56
timestamp 1666464484
transform 1 0 56674 0 1 69427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_57
timestamp 1666464484
transform 1 0 56674 0 1 71227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_58
timestamp 1666464484
transform 1 0 56674 0 1 73027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_59
timestamp 1666464484
transform 1 0 56674 0 1 74827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_60
timestamp 1666464484
transform 1 0 56674 0 1 76627
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_61
timestamp 1666464484
transform 1 0 56674 0 1 78427
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_62
timestamp 1666464484
transform 1 0 56674 0 1 80227
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_63
timestamp 1666464484
transform 1 0 56674 0 1 82027
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_64
timestamp 1666464484
transform 1 0 56674 0 1 83827
box 0 0 1 1
use M2_M1$$199747628_512x8m81  M2_M1$$199747628_512x8m81_65
timestamp 1666464484
transform 1 0 56674 0 1 85627
box 0 0 1 1
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_512x8m81  M2_M1$$201260076_512x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_512x8m81  M2_M1$$201261100_512x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 4126
box -170 -502 170 502
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1666464484
transform 1 0 62228 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1666464484
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1666464484
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_3
timestamp 1666464484
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_4
timestamp 1666464484
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_5
timestamp 1666464484
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_6
timestamp 1666464484
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_7
timestamp 1666464484
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_8
timestamp 1666464484
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_9
timestamp 1666464484
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_10
timestamp 1666464484
transform 1 0 40701 0 1 3256
box 0 0 1 1
use M2_M1431059130203_512x8m81  M2_M1431059130203_512x8m81_0
timestamp 1666464484
transform 1 0 25662 0 1 34778
box -286 -224 286 224
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_0
timestamp 1666464484
transform 1 0 25662 0 1 94623
box -286 -162 286 162
use M2_M1431059130204_512x8m81  M2_M1431059130204_512x8m81_1
timestamp 1666464484
transform 1 0 59141 0 1 94623
box -286 -162 286 162
use M2_M1431059130208_512x8m81  M2_M1431059130208_512x8m81_0
timestamp 1666464484
transform 1 0 60601 0 1 35416
box 0 0 1 1
use M2_M14310591302012_512x8m81  M2_M14310591302012_512x8m81_0
timestamp 1666464484
transform 1 0 27599 0 1 34778
box -162 -224 162 224
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 12783
box -170 -1046 170 1046
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 15671
box -170 -1046 170 1046
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 15463
box -170 -1046 170 1046
use M3_M2$$201248812_512x8m81  M3_M2$$201248812_512x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 13112
box -170 -1046 170 1046
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 10834
box -170 -611 170 611
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 8835
box -170 -611 170 611
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 10834
box -170 -611 170 611
use M3_M2$$201249836_512x8m81  M3_M2$$201249836_512x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 8835
box -170 -611 170 611
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_0
timestamp 1666464484
transform -1 0 56505 0 1 6590
box -381 -284 381 284
use M3_M2$$201250860_512x8m81  M3_M2$$201250860_512x8m81_1
timestamp 1666464484
transform 1 0 28618 0 1 6590
box -381 -284 381 284
use M3_M2$$201251884_512x8m81  M3_M2$$201251884_512x8m81_0
timestamp 1666464484
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_512x8m81  M3_M2$$201252908_512x8m81_0
timestamp 1666464484
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201253932_512x8m81  M3_M2$$201253932_512x8m81_0
timestamp 1666464484
transform 1 0 57515 0 1 8162
box -170 -1155 170 730
use M3_M2$$201254956_512x8m81  M3_M2$$201254956_512x8m81_0
timestamp 1666464484
transform 1 0 27608 0 1 13768
box -170 -502 170 502
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_0
timestamp 1666464484
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_1
timestamp 1666464484
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_2
timestamp 1666464484
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_3
timestamp 1666464484
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_4
timestamp 1666464484
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_5
timestamp 1666464484
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_6
timestamp 1666464484
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_7
timestamp 1666464484
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_8
timestamp 1666464484
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_9
timestamp 1666464484
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_10
timestamp 1666464484
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_11
timestamp 1666464484
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_12
timestamp 1666464484
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_13
timestamp 1666464484
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_14
timestamp 1666464484
transform 1 0 28449 0 1 82027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_15
timestamp 1666464484
transform 1 0 28449 0 1 80227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_16
timestamp 1666464484
transform 1 0 28449 0 1 78427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_17
timestamp 1666464484
transform 1 0 28449 0 1 76627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_18
timestamp 1666464484
transform 1 0 28449 0 1 74827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_19
timestamp 1666464484
transform 1 0 28449 0 1 73027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_20
timestamp 1666464484
transform 1 0 28449 0 1 71227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_21
timestamp 1666464484
transform 1 0 28449 0 1 69427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_22
timestamp 1666464484
transform 1 0 28449 0 1 67627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_23
timestamp 1666464484
transform 1 0 28449 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_24
timestamp 1666464484
transform 1 0 28449 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_25
timestamp 1666464484
transform 1 0 28449 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_26
timestamp 1666464484
transform 1 0 28449 0 1 60427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_27
timestamp 1666464484
transform 1 0 28449 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_28
timestamp 1666464484
transform 1 0 28449 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_29
timestamp 1666464484
transform 1 0 28449 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_30
timestamp 1666464484
transform 1 0 28449 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_31
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_32
timestamp 1666464484
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_33
timestamp 1666464484
transform 1 0 28449 0 1 94627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_34
timestamp 1666464484
transform 1 0 28449 0 1 92827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_35
timestamp 1666464484
transform 1 0 28449 0 1 91027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_36
timestamp 1666464484
transform 1 0 28449 0 1 89227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_37
timestamp 1666464484
transform 1 0 28449 0 1 87427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_38
timestamp 1666464484
transform 1 0 28449 0 1 85627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_39
timestamp 1666464484
transform 1 0 28449 0 1 83827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_40
timestamp 1666464484
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_41
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_42
timestamp 1666464484
transform 1 0 56674 0 1 53227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_43
timestamp 1666464484
transform 1 0 56674 0 1 55027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_44
timestamp 1666464484
transform 1 0 56674 0 1 56827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_45
timestamp 1666464484
transform 1 0 56674 0 1 58627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_46
timestamp 1666464484
transform 1 0 56674 0 1 60427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_47
timestamp 1666464484
transform 1 0 56674 0 1 62227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_48
timestamp 1666464484
transform 1 0 56674 0 1 64027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_49
timestamp 1666464484
transform 1 0 56674 0 1 65827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_50
timestamp 1666464484
transform 1 0 56674 0 1 67627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_51
timestamp 1666464484
transform 1 0 56674 0 1 69427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_52
timestamp 1666464484
transform 1 0 56674 0 1 71227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_53
timestamp 1666464484
transform 1 0 56674 0 1 73027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_54
timestamp 1666464484
transform 1 0 56674 0 1 74827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_55
timestamp 1666464484
transform 1 0 56674 0 1 76627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_56
timestamp 1666464484
transform 1 0 56674 0 1 78427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_57
timestamp 1666464484
transform 1 0 56674 0 1 80227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_58
timestamp 1666464484
transform 1 0 56674 0 1 82027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_59
timestamp 1666464484
transform 1 0 56674 0 1 83827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_60
timestamp 1666464484
transform 1 0 56674 0 1 85627
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_61
timestamp 1666464484
transform 1 0 56674 0 1 87427
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_62
timestamp 1666464484
transform 1 0 56674 0 1 89227
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_63
timestamp 1666464484
transform 1 0 56674 0 1 91027
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_64
timestamp 1666464484
transform 1 0 56674 0 1 92827
box 0 0 1 1
use M3_M2$$201258028_512x8m81  M3_M2$$201258028_512x8m81_65
timestamp 1666464484
transform 1 0 56674 0 1 94627
box 0 0 1 1
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 30897
box -170 -393 170 393
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 32786
box -170 -393 170 393
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 32786
box -170 -393 170 393
use M3_M2$$201412652_512x8m81  M3_M2$$201412652_512x8m81_3
timestamp 1666464484
transform 1 0 27608 0 1 30897
box -170 -393 170 393
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_1
timestamp 1666464484
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_512x8m81  M3_M2$$201413676_512x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 33221
box -170 -828 170 828
use M3_M2$$201414700_512x8m81  M3_M2$$201414700_512x8m81_1
timestamp 1666464484
transform 1 0 26993 0 1 33221
box -170 -828 170 828
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 28743
box -170 -1264 170 1264
use M3_M2$$201415724_512x8m81  M3_M2$$201415724_512x8m81_1
timestamp 1666464484
transform 1 0 26993 0 1 28743
box -170 -1264 170 1264
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_2
timestamp 1666464484
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_3
timestamp 1666464484
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_4
timestamp 1666464484
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_5
timestamp 1666464484
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_6
timestamp 1666464484
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_7
timestamp 1666464484
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_8
timestamp 1666464484
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_9
timestamp 1666464484
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_512x8m81  M3_M2$$201416748_512x8m81_10
timestamp 1666464484
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_0
timestamp 1666464484
transform 0 -1 49977 1 0 8925
box 0 0 1 1
use M3_M2431059130201_512x8m81  M3_M2431059130201_512x8m81_1
timestamp 1666464484
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431059130202_512x8m81  M3_M2431059130202_512x8m81_0
timestamp 1666464484
transform 1 0 25662 0 1 34778
box -286 -224 286 224
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_0
timestamp 1666464484
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_1
timestamp 1666464484
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_2
timestamp 1666464484
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_3
timestamp 1666464484
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_4
timestamp 1666464484
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_5
timestamp 1666464484
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_6
timestamp 1666464484
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_7
timestamp 1666464484
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_8
timestamp 1666464484
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_9
timestamp 1666464484
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_10
timestamp 1666464484
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_11
timestamp 1666464484
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_12
timestamp 1666464484
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_13
timestamp 1666464484
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_14
timestamp 1666464484
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_15
timestamp 1666464484
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_16
timestamp 1666464484
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_17
timestamp 1666464484
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_18
timestamp 1666464484
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431059130205_512x8m81  M3_M2431059130205_512x8m81_19
timestamp 1666464484
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431059130206_512x8m81  M3_M2431059130206_512x8m81_0
timestamp 1666464484
transform 1 0 27599 0 1 34778
box -162 -224 162 224
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1666464484
transform 1 0 43880 0 1 3022
box 0 0 1 1
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_0
timestamp 1666464484
transform 1 0 59149 0 1 31146
box -286 -162 286 162
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_1
timestamp 1666464484
transform 1 0 59149 0 1 30701
box -286 -162 286 162
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_2
timestamp 1666464484
transform 1 0 25674 0 1 31096
box -286 -162 286 162
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_3
timestamp 1666464484
transform 1 0 25674 0 1 30641
box -286 -162 286 162
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_4
timestamp 1666464484
transform 1 0 25662 0 1 94623
box -286 -162 286 162
use M3_M2431059130209_512x8m81  M3_M2431059130209_512x8m81_5
timestamp 1666464484
transform 1 0 59141 0 1 94623
box -286 -162 286 162
use M3_M24310591302011_512x8m81  M3_M24310591302011_512x8m81_0
timestamp 1666464484
transform 1 0 59154 0 1 34778
box -348 -224 348 224
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_0
timestamp 1666464484
transform 1 0 58126 0 1 23631
box -142 -454 142 454
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_1
timestamp 1666464484
transform 1 0 57495 0 1 22479
box -142 -454 142 454
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_2
timestamp 1666464484
transform 1 0 26990 0 1 23631
box -142 -454 142 454
use M3_M24310591302013_512x8m81  M3_M24310591302013_512x8m81_3
timestamp 1666464484
transform 1 0 27607 0 1 22492
box -142 -454 142 454
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_0
timestamp 1666464484
transform 1 0 59135 0 1 27399
box -286 -906 286 906
use M3_M24310591302015_512x8m81  M3_M24310591302015_512x8m81_1
timestamp 1666464484
transform 1 0 25680 0 1 27421
box -286 -906 286 906
use control_512x8_512x8m81  control_512x8_512x8m81_0
timestamp 1666464484
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use lcol4_512_512x8m81  lcol4_512_512x8m81_0
timestamp 1666464484
transform 1 0 2921 0 1 5019
box -1235 -3416 22810 89707
use m2m3_512x8m81  m2m3_512x8m81_0
timestamp 1666464484
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use power_a_512x8m81  power_a_512x8m81_0
timestamp 1666464484
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_1
timestamp 1666464484
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_2
timestamp 1666464484
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_3
timestamp 1666464484
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_4
timestamp 1666464484
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_5
timestamp 1666464484
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_6
timestamp 1666464484
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_7
timestamp 1666464484
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_8
timestamp 1666464484
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_9
timestamp 1666464484
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_10
timestamp 1666464484
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_11
timestamp 1666464484
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_12
timestamp 1666464484
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_13
timestamp 1666464484
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_14
timestamp 1666464484
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_15
timestamp 1666464484
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_a_512x8m81  power_a_512x8m81_16
timestamp 1666464484
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_0
timestamp 1666464484
transform 1 0 15448 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_1
timestamp 1666464484
transform 1 0 10048 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_2
timestamp 1666464484
transform 1 0 4648 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_3
timestamp 1666464484
transform 1 0 75024 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_4
timestamp 1666464484
transform 1 0 69624 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_5
timestamp 1666464484
transform 1 0 64224 0 1 94546
box -511 630 1714 2430
use power_route_01_a_512x8m81  power_route_01_a_512x8m81_6
timestamp 1666464484
transform 1 0 46824 0 1 94546
box -511 630 1714 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_0
timestamp 1666464484
transform -1 0 41719 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_1
timestamp 1666464484
transform -1 0 39074 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_2
timestamp 1666464484
transform -1 0 35904 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_3
timestamp 1666464484
transform -1 0 31199 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_4
timestamp 1666464484
transform -1 0 27061 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_5
timestamp 1666464484
transform -1 0 21142 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_6
timestamp 1666464484
transform -1 0 80718 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_7
timestamp 1666464484
transform -1 0 58036 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_8
timestamp 1666464484
transform -1 0 85155 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_9
timestamp 1666464484
transform -1 0 54751 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_10
timestamp 1666464484
transform -1 0 49390 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_11
timestamp 1666464484
transform -1 0 45558 0 1 94546
box -511 630 489 2430
use power_route_01_b_512x8m81  power_route_01_b_512x8m81_12
timestamp 1666464484
transform -1 0 53058 0 1 94546
box -511 630 489 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_0
timestamp 1666464484
transform -1 0 26872 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_1
timestamp 1666464484
transform -1 0 41596 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_2
timestamp 1666464484
transform -1 0 38662 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_3
timestamp 1666464484
transform -1 0 35738 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_4
timestamp 1666464484
transform -1 0 34095 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_5
timestamp 1666464484
transform -1 0 30987 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_6
timestamp 1666464484
transform -1 0 29591 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_7
timestamp 1666464484
transform -1 0 60505 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_8
timestamp 1666464484
transform -1 0 52179 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_9
timestamp 1666464484
transform -1 0 45427 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_10
timestamp 1666464484
transform -1 0 57704 0 1 94546
box 714 1822 1714 2430
use power_route_01_c_512x8m81  power_route_01_c_512x8m81_11
timestamp 1666464484
transform -1 0 44144 0 1 94546
box 714 1822 1714 2430
use power_route_512x8m81  power_route_512x8m81_0
timestamp 1666464484
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 99039
use rcol4_512_512x8m81  rcol4_512_512x8m81_0
timestamp 1666464484
transform 1 0 60511 0 1 5019
box -1090 -3398 24835 89717
use xdec64_512x8m81  xdec64_512x8m81_0
timestamp 1666464484
transform 1 0 28677 0 1 36127
box -3364 -228 31133 58748
<< labels >>
flabel metal3 s 0 93376 1706 94076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 91576 1706 92276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 89776 1706 90476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87976 1706 88676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 86176 1706 86876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 2626 96368 3626 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 5362 96368 6362 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 8026 96368 9026 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 10762 96368 11762 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 13426 96368 14426 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 84376 1706 85076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 82576 1706 83276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 80776 1706 81476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 78976 1706 79676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 77176 1706 77876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 75376 1706 76076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 73576 1706 74276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 71776 1706 72476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 16162 96368 17162 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 18826 96368 19826 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 22258 96368 23258 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 25158 96368 26158 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 26435 3011 28416 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 6921 26434 8163 28412 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 69976 1706 70676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 68176 1706 68876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 66376 1706 67076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 64576 1706 65276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 62776 1706 63476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17721 26434 18963 28412 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 60976 1706 61676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 26435 26070 28412 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 59176 1706 59876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23425 26434 27828 26890 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 34536 1014 35326 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 35126 24917 35326 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 34536 27830 35016 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 27877 96368 28877 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 57376 1706 58076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 55576 1706 56276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 53776 1706 54476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 51976 1706 52676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 50176 1706 50876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 48376 1706 49076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 46576 1706 47276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 44776 1706 45476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29273 96368 30273 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 32381 96368 33381 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 34024 96368 35024 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8152 1014 9515 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8152 3011 9514 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 36948 96368 37948 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 39882 96368 40882 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 42430 96368 43430 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 43713 96368 44713 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 47538 96368 48538 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2226 8154 28729 9515 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 8153 24250 9514 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 1401 95176 2401 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 4137 95176 5137 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 6801 95176 7801 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 9537 95176 10537 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50465 96368 51465 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 12201 95176 13201 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 55990 96368 56990 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58791 96368 59791 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 62202 96368 63202 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 14937 95176 15937 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 17601 95176 18601 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 20653 95176 21653 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23483 95176 24483 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26572 95176 27572 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30710 95176 31710 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 35415 95176 36415 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 38585 95176 39585 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 41230 95176 42230 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 64938 96368 65938 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 67602 96368 68602 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 70338 96368 71338 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 73002 96368 74002 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 75738 96368 76738 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 78402 96368 79402 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 45069 95176 46069 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 46313 95176 47313 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 48901 95176 49901 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 52569 95176 53569 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 81834 96368 82834 96976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94276 1014 94976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 25376 94461 25948 94785 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94476 27272 94776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30402 94526 54622 94728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 94527 86372 94728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58855 94461 59427 94785 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 58855 94476 86372 94776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 94276 86372 94976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 54262 95176 55262 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57547 95176 58547 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92476 1014 93176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 60977 95176 61977 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92676 27272 92976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 63713 95176 64713 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 66377 95176 67377 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 69113 95176 70113 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 71777 95176 72777 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 74513 95176 75513 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 77177 95176 78177 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 80229 95176 81229 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83059 95176 84059 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 92726 54622 92928 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 95176 85666 96976 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 92727 86372 92928 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 95176 86372 96176 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 92676 86372 92976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 93376 86372 94076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 92476 86372 93176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 91576 86372 92276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 90676 1014 91376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 90876 27272 91176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 90926 54622 91128 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 90927 86372 91128 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 90876 86372 91176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 90676 86372 91376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 88876 1014 89576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 89776 86372 90476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 87976 86372 88676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 86176 86372 86876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 89076 27272 89376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 89126 54622 89328 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 89127 86372 89328 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 89076 86372 89376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 84376 86372 85076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 82576 86372 83276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 80776 86372 81476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 78976 86372 79676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 77176 86372 77876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 75376 86372 76076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 73576 86372 74276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 71776 86372 72476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 69976 86372 70676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 68176 86372 68876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 66376 86372 67076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 64576 86372 65276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 62776 86372 63476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 88876 86372 89576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 60976 86372 61676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87076 1014 87776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 87276 27272 87576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 59176 86372 59876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 57376 86372 58076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 55576 86372 56276 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 53776 86372 54476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 51976 86372 52676 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 50176 86372 50876 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 48376 86372 49076 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 46576 86372 47276 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 87326 54622 87528 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 44776 86372 45476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 87327 86372 87528 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 87276 86372 87576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 87076 86372 87776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 85276 1014 85976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 85476 27272 85776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 85526 54622 85728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 85527 86372 85728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 85476 86372 85776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 85276 86372 85976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 83476 1014 84176 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 83676 27272 83976 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 83726 54622 83928 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 83727 86372 83928 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 59421 83676 86372 83976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 83476 86372 84176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 81676 1014 82376 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 81876 27272 82176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 81926 54622 82128 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 81927 86372 82128 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 81876 86372 82176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 81676 86372 82376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 79876 1014 80576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 80076 27272 80376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 30403 80126 54622 80328 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 80127 86372 80328 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61825 18015 83763 20739 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61807 18016 86372 20739 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 34741 9972 41516 12570 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29478 10756 41516 12570 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12570 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 26772 11844 58351 12570 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 61773 13461 86372 14177 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 80076 86372 80376 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 79876 86372 80576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78076 1014 78776 0 FreeSans 2000 180 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78276 27272 78576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 26772 12035 84999 12570 0 FreeSans 2000 180 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 78326 54622 78528 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 78327 86372 78528 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 78276 86372 78576 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 61802 8153 86372 9514 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 85358 78076 86372 78776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76276 1014 76976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 57909 8154 72434 9515 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76476 27272 76776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 72602 8152 83234 9515 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 76526 54622 76728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 61825 8152 86372 9514 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 76527 86372 76728 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 8152 86372 9515 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 59421 76476 86372 76776 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 85358 76276 86372 76976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 4060 1712 5629 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 74476 1014 75176 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 5173 3011 5629 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 0 74676 27272 74976 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
flabel metal3 s 0 5174 24250 5629 0 FreeSans 2000 0 0 0 VDD
port 29 nsew power bidirectional
flabel metal3 s 30403 74726 54622 74928 0 FreeSans 2000 0 0 0 VSS
port 30 nsew ground bidirectional
rlabel metal2 s 27936 0 28160 200 4 CLK
port 11 nsew signal input
rlabel metal2 s 1864 0 2088 200 4 D[0]
port 19 nsew signal input
rlabel metal2 s 29006 0 29230 200 4 A[8]
port 1 nsew signal input
rlabel metal2 s 29705 0 29929 200 4 A[7]
port 2 nsew signal input
rlabel metal2 s 30859 0 31083 200 4 A[2]
port 7 nsew signal input
rlabel metal2 s 32552 0 32776 200 4 A[1]
port 8 nsew signal input
rlabel metal2 s 34243 0 34467 200 4 A[0]
port 9 nsew signal input
rlabel metal2 s 14127 0 14351 200 4 Q[2]
port 26 nsew signal output
rlabel metal2 s 22279 0 22503 200 4 Q[3]
port 25 nsew signal output
rlabel metal2 s 50342 0 50566 200 4 CEN
port 10 nsew signal input
rlabel metal2 s 54417 0 54641 200 4 A[5]
port 4 nsew signal input
rlabel metal2 s 53772 0 53996 200 4 A[6]
port 3 nsew signal input
rlabel metal2 s 55164 0 55388 200 4 A[4]
port 5 nsew signal input
rlabel metal2 s 23404 0 23628 200 4 WEN[3]
port 35 nsew signal input
rlabel metal2 s 83372 0 83596 200 4 D[7]
port 12 nsew signal input
rlabel metal2 s 81855 0 82079 200 4 Q[7]
port 21 nsew signal output
rlabel metal2 s 23795 0 24019 200 4 D[3]
port 16 nsew signal input
rlabel metal2 s 12206 0 12430 200 4 D[1]
port 18 nsew signal input
rlabel metal2 s 13454 0 13678 200 4 D[2]
port 17 nsew signal input
rlabel metal2 s 56265 0 56489 200 4 A[3]
port 6 nsew signal input
rlabel metal2 s 11533 0 11757 200 4 Q[1]
port 27 nsew signal output
rlabel metal2 s 73703 0 73927 200 4 Q[6]
port 22 nsew signal output
rlabel metal2 s 71782 0 72006 200 4 D[5]
port 14 nsew signal input
rlabel metal2 s 62958 0 63182 200 4 Q[4]
port 24 nsew signal output
rlabel metal2 s 72180 0 72404 200 4 WEN[5]
port 33 nsew signal input
rlabel metal2 s 13054 0 13278 200 4 WEN[2]
port 36 nsew signal input
rlabel metal2 s 12604 0 12828 200 4 WEN[1]
port 37 nsew signal input
rlabel metal2 s 62115 0 62339 200 4 WEN[4]
port 34 nsew signal input
rlabel metal2 s 82695 0 82919 200 4 WEN[7]
port 31 nsew signal input
rlabel metal2 s 72630 0 72854 200 4 WEN[6]
port 32 nsew signal input
rlabel metal2 s 61447 0 61671 200 4 D[4]
port 15 nsew signal input
rlabel metal2 s 73030 0 73254 200 4 D[6]
port 13 nsew signal input
rlabel metal2 s 71109 0 71333 200 4 Q[5]
port 23 nsew signal output
rlabel metal2 s 3380 0 3604 200 4 Q[0]
port 28 nsew signal output
rlabel metal2 s 40588 0 40812 200 4 GWEN
port 20 nsew signal input
rlabel metal2 s 2539 0 2763 200 4 WEN[0]
port 38 nsew signal input
flabel space 0 200 0 200 3 FreeSans 2000 0 0 0 & Metric 1.00
flabel space 0 600 0 600 3 FreeSans 2000 0 0 0 & Version 2015q2v1
flabel space 0 1000 0 1000 3 FreeSans 2000 0 0 0 & Product GF018_5VGreen_SRAM_1P_512x8M8WM1
flabel metal3 0 1400 0 1400 3 FreeSans 2000 0 0 0 & Vendor GLOBALFOUNDRIES
rlabel metal3 s 0 4060 24341 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 29 nsew power bidirectional
rlabel metal3 s 0 74727 86372 74928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 74676 86372 74976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 74476 86372 75176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72676 1014 73376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72876 27272 73176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 72926 54622 73128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 72927 86372 73128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 72876 86372 73176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 72676 86372 73376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 70876 1014 71576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71076 27272 71376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 71126 54622 71328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 71127 86372 71328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 71076 86372 71376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 70876 86372 71576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69076 1014 69776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69276 27272 69576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 69326 54622 69528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 69327 86372 69528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 69276 86372 69576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 69076 86372 69776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67276 1014 67976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67476 27272 67776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 67526 54622 67728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 67527 86372 67728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 67476 86372 67776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 67276 86372 67976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65476 1014 66176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65676 27272 65976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 65726 54622 65928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 65727 86372 65928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 65676 86372 65976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 65476 86372 66176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63676 1014 64376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63876 27272 64176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 63926 54622 64128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 63927 86372 64128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 63876 86372 64176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 63676 86372 64376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 61876 1014 62576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62076 27272 62376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 62126 54622 62328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 62127 86372 62328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 62076 86372 62376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 61876 86372 62576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60076 1014 60776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60276 27272 60576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 60326 54622 60528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 60327 86372 60528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 60276 86372 60576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 60076 86372 60776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58276 1014 58976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58476 27272 58776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 58526 54622 58728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 58527 86372 58728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 58476 86372 58776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 58276 86372 58976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56476 1014 57176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56676 27272 56976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 56726 54622 56928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 56727 86372 56928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 56676 86372 56976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 56476 86372 57176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54676 1014 55376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54876 27272 55176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 54926 54622 55128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 54927 86372 55128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 54876 86372 55176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 54676 86372 55376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 52876 1014 53576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53076 27272 53376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 53126 54622 53328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 53127 86372 53328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 53076 86372 53376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 52876 86372 53576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51076 1014 51776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51276 27272 51576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 51326 54622 51528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 51327 86372 51528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 51276 86372 51576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 51076 86372 51776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49276 1014 49976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49476 27272 49776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 49526 54622 49728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 49527 86372 49728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 49476 86372 49776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 49276 86372 49976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47476 1014 48176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47676 27272 47976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 47726 54622 47928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 47727 86372 47928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 47676 86372 47976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 47476 86372 48176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45676 1014 46376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45876 27272 46176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 45926 54622 46128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 45927 86372 46128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 45876 86372 46176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 45676 86372 46376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 43876 1014 44576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44076 27272 44376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 44127 86372 44328 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 42327 86372 42528 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 40527 86372 40728 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 38727 86372 38928 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 36927 86372 37128 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60460 35158 86372 35298 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58791 34536 86372 35016 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 34536 86372 35326 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83360 35126 86372 35326 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28412 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 26435 86372 28416 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 57681 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 22291 57681 23199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42261 10740 86372 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8930 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 1014 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 1 VSS
port 30 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 30 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 96976
string GDS_END 2941440
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2876172
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 232.665 4.660 232.665 0.000 
<< end >>
