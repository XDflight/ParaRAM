magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 3136 844
rect 69 496 115 724
rect 468 430 550 674
rect 1249 569 1317 724
rect 58 354 318 430
rect 373 354 550 430
rect 1938 584 1984 724
rect 262 60 330 199
rect 1213 60 1281 215
rect 2327 492 2373 724
rect 2740 580 2786 724
rect 2832 466 3046 654
rect 2043 318 2213 353
rect 2043 307 2551 318
rect 2157 242 2551 307
rect 1964 60 2010 169
rect 2956 224 3046 466
rect 2740 60 2786 161
rect 2940 112 3046 224
rect 0 -60 3136 60
<< obsm1 >>
rect 762 512 808 625
rect 1464 632 1879 678
rect 600 466 1087 512
rect 38 245 423 292
rect 38 153 106 245
rect 377 199 423 245
rect 600 199 646 466
rect 692 374 987 420
rect 692 289 738 374
rect 1041 315 1087 466
rect 1464 407 1510 632
rect 1729 407 1786 570
rect 1833 538 1879 632
rect 2040 632 2281 678
rect 2040 538 2086 632
rect 1833 491 2086 538
rect 2143 445 2189 570
rect 1137 361 1510 407
rect 1041 268 1416 315
rect 377 153 554 199
rect 600 153 778 199
rect 1464 156 1510 361
rect 1583 361 1786 407
rect 1849 399 2189 445
rect 2235 445 2281 632
rect 2536 534 2582 650
rect 2536 488 2775 534
rect 2235 442 2453 445
rect 2235 399 2683 442
rect 1583 152 1655 361
rect 1849 261 1897 399
rect 2402 393 2683 399
rect 2729 405 2775 488
rect 2729 337 2910 405
rect 2729 307 2775 337
rect 1849 215 2102 261
rect 2602 253 2775 307
rect 1583 106 1815 152
rect 2056 152 2102 215
rect 2602 152 2648 253
rect 2056 106 2247 152
rect 2319 106 2648 152
<< labels >>
rlabel metal1 s 2043 318 2213 353 6 CLK
port 1 nsew clock input
rlabel metal1 s 2043 307 2551 318 6 CLK
port 1 nsew clock input
rlabel metal1 s 2157 242 2551 307 6 CLK
port 1 nsew clock input
rlabel metal1 s 468 430 550 674 6 E
port 2 nsew default input
rlabel metal1 s 373 354 550 430 6 E
port 2 nsew default input
rlabel metal1 s 58 354 318 430 6 TE
port 3 nsew default input
rlabel metal1 s 2832 466 3046 654 6 Q
port 4 nsew default output
rlabel metal1 s 2956 224 3046 466 6 Q
port 4 nsew default output
rlabel metal1 s 2940 112 3046 224 6 Q
port 4 nsew default output
rlabel metal1 s 0 724 3136 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 584 2786 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 584 2373 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1938 584 1984 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 584 1317 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 584 115 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2740 580 2786 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 580 2373 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 580 1317 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 580 115 584 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 569 2373 580 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1249 569 1317 580 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 569 115 580 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 496 2373 569 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 69 496 115 569 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2327 492 2373 496 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1213 199 1281 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 169 1281 199 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 169 330 199 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1964 161 2010 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 161 1281 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 161 330 169 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2740 60 2786 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1964 60 2010 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1213 60 1281 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 3136 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3136 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 449430
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 442292
<< end >>
