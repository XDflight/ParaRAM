magic
tech gf180mcuA
timestamp 1666464484
<< metal1 >>
rect 0 147 44 159
rect 11 106 16 147
rect 28 45 33 46
rect 26 39 36 45
rect 11 9 16 33
rect 28 16 33 39
rect 0 -3 44 9
<< obsm1 >>
rect 28 99 33 140
rect 23 94 33 99
<< metal2 >>
rect 10 154 18 155
rect 9 148 19 154
rect 10 147 18 148
rect 26 38 36 46
rect 10 8 18 9
rect 9 2 19 8
rect 10 1 18 2
<< labels >>
rlabel metal2 s 10 147 18 155 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 147 44 159 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 2 nsew ground bidirectional
rlabel metal1 s 11 -3 16 33 6 VSS
port 2 nsew ground bidirectional
rlabel metal1 s 0 -3 44 9 6 VSS
port 2 nsew ground bidirectional
rlabel metal2 s 26 38 36 46 6 Y
port 3 nsew signal output
rlabel metal1 s 28 16 33 46 6 Y
port 3 nsew signal output
rlabel metal1 s 26 39 36 45 6 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 44 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
