magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 4032 844
rect 262 586 330 724
rect 648 569 716 724
rect 1535 689 1603 724
rect 56 353 318 426
rect 578 354 806 430
rect 262 60 330 210
rect 630 60 698 215
rect 2055 601 2123 724
rect 2859 601 2927 724
rect 1491 60 1559 215
rect 3342 506 3388 724
rect 2818 354 3057 430
rect 3690 506 3736 724
rect 3809 438 3963 676
rect 3311 60 3379 210
rect 3885 232 3963 438
rect 3690 60 3736 153
rect 3860 110 3963 232
rect 0 -60 4032 60
<< obsm1 >>
rect 69 519 115 645
rect 477 523 523 645
rect 762 632 1023 678
rect 1654 643 1983 678
rect 762 523 808 632
rect 69 472 418 519
rect 372 302 418 472
rect 49 256 418 302
rect 477 476 808 523
rect 49 162 95 256
rect 477 230 524 476
rect 477 162 543 230
rect 854 158 922 586
rect 977 386 1023 632
rect 1223 632 1983 643
rect 1223 597 1700 632
rect 1069 399 1115 597
rect 1223 448 1291 597
rect 1807 491 1875 586
rect 1937 555 1983 632
rect 2169 613 2463 659
rect 2169 555 2215 613
rect 1937 508 2215 555
rect 1403 462 1875 491
rect 2261 462 2329 556
rect 1403 445 2329 462
rect 1807 416 2329 445
rect 2386 510 2579 556
rect 2726 555 2772 569
rect 3074 555 3120 577
rect 1069 353 1647 399
rect 1069 158 1135 353
rect 1200 261 1668 307
rect 1622 152 1668 261
rect 1975 198 2043 416
rect 2162 152 2208 323
rect 2386 226 2432 510
rect 2726 508 3120 555
rect 2726 244 2772 508
rect 3546 421 3592 676
rect 3151 372 3592 421
rect 3546 368 3592 372
rect 3176 279 3467 326
rect 3546 300 3824 368
rect 2254 158 2432 226
rect 2511 198 2899 244
rect 1622 106 2208 152
rect 2386 152 2432 158
rect 3176 152 3222 279
rect 2386 106 3222 152
rect 3546 161 3592 300
<< labels >>
rlabel metal1 s 578 354 806 430 6 D
port 1 nsew default input
rlabel metal1 s 2818 354 3057 430 6 SETN
port 2 nsew default input
rlabel metal1 s 56 353 318 426 6 CLK
port 3 nsew clock input
rlabel metal1 s 3809 438 3963 676 6 Q
port 4 nsew default output
rlabel metal1 s 3885 232 3963 438 6 Q
port 4 nsew default output
rlabel metal1 s 3860 110 3963 232 6 Q
port 4 nsew default output
rlabel metal1 s 0 724 4032 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3690 689 3736 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3342 689 3388 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2859 689 2927 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2055 689 2123 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1535 689 1603 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 689 716 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 689 330 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3690 601 3736 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3342 601 3388 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2859 601 2927 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2055 601 2123 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 601 716 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 601 330 689 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3690 586 3736 601 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3342 586 3388 601 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 586 716 601 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 262 586 330 601 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3690 569 3736 586 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3342 569 3388 586 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 648 569 716 586 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3690 506 3736 569 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3342 506 3388 569 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1491 210 1559 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 630 210 698 215 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3311 153 3379 210 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1491 153 1559 210 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 630 153 698 210 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 153 330 210 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3690 60 3736 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3311 60 3379 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1491 60 1559 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 630 60 698 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 60 330 153 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4032 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1038160
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1029548
<< end >>
