magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -68 622 668 968
<< pwell >>
rect -68 -68 668 622
<< mvnmos >>
rect 126 342 246 532
rect 354 342 474 532
rect 36 52 156 206
rect 444 52 564 206
<< mvpmos >>
rect 126 712 246 832
rect 354 712 474 832
<< mvndiff >>
rect 36 413 126 532
rect 36 367 49 413
rect 95 367 126 413
rect 36 342 126 367
rect 246 342 354 532
rect 474 413 564 532
rect 474 367 505 413
rect 551 367 564 413
rect 474 342 564 367
rect 36 270 96 342
rect 270 331 330 342
rect 270 285 277 331
rect 323 285 330 331
rect 36 206 156 270
rect 270 266 330 285
rect 504 270 564 342
rect 444 206 564 270
rect 36 23 156 52
rect 36 -23 73 23
rect 119 -23 156 23
rect 36 -42 156 -23
rect 444 23 564 52
rect 444 -23 481 23
rect 527 -23 564 23
rect 444 -42 564 -23
<< mvpdiff >>
rect 270 923 330 942
rect 270 877 277 923
rect 323 877 330 923
rect 270 832 330 877
rect 36 771 126 832
rect 36 725 49 771
rect 95 725 126 771
rect 36 712 126 725
rect 246 712 354 832
rect 474 771 564 832
rect 474 725 505 771
rect 551 725 564 771
rect 474 712 564 725
<< mvndiffc >>
rect 49 367 95 413
rect 505 367 551 413
rect 277 285 323 331
rect 73 -23 119 23
rect 481 -23 527 23
<< mvpdiffc >>
rect 277 877 323 923
rect 49 725 95 771
rect 505 725 551 771
<< polysilicon >>
rect 126 832 246 876
rect 354 832 474 876
rect 126 631 246 712
rect 126 585 187 631
rect 233 585 246 631
rect 126 532 246 585
rect 354 659 474 712
rect 354 613 367 659
rect 413 613 474 659
rect 354 532 474 613
rect 126 298 246 342
rect 354 298 474 342
rect -36 52 36 206
rect 156 52 444 206
rect 564 52 636 206
<< polycontact >>
rect 187 585 233 631
rect 367 613 413 659
<< metal1 >>
rect -36 923 636 950
rect -36 877 277 923
rect 323 877 636 923
rect -36 850 636 877
rect 38 771 414 790
rect 38 725 49 771
rect 95 725 414 771
rect 38 716 414 725
rect 38 413 112 716
rect 340 659 414 716
rect 186 631 260 650
rect 186 585 187 631
rect 233 585 260 631
rect 340 613 367 659
rect 413 613 414 659
rect 340 594 414 613
rect 488 771 562 790
rect 488 725 505 771
rect 551 725 562 771
rect 186 528 260 585
rect 488 528 562 725
rect 186 454 562 528
rect 38 367 49 413
rect 95 367 112 413
rect 488 413 562 454
rect 38 348 112 367
rect 248 331 352 374
rect 488 367 505 413
rect 551 367 562 413
rect 488 348 562 367
rect 248 285 277 331
rect 323 285 352 331
rect 248 258 352 285
rect -36 138 636 258
rect 36 23 248 50
rect 36 -23 73 23
rect 119 -23 248 23
rect 36 -50 248 -23
rect 352 23 564 50
rect 352 -23 481 23
rect 527 -23 564 23
rect 352 -50 564 -23
<< metal2 >>
rect 90 -50 210 950
rect 390 -50 510 950
<< metal3 >>
rect -36 330 636 690
<< properties >>
string FIXED_BBOX -68 -68 668 968
string GDS_END 409020
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 406664
<< end >>
