magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 120
rect 224 0 344 120
<< mvndiff >>
rect -88 83 0 120
rect -88 37 -75 83
rect -29 37 0 83
rect -88 0 0 37
rect 120 83 224 120
rect 120 37 149 83
rect 195 37 224 83
rect 120 0 224 37
rect 344 83 432 120
rect 344 37 373 83
rect 419 37 432 83
rect 344 0 432 37
<< mvndiffc >>
rect -75 37 -29 83
rect 149 37 195 83
rect 373 37 419 83
<< polysilicon >>
rect 0 120 120 164
rect 224 120 344 164
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 83 -29 120
rect -75 0 -29 37
rect 149 83 195 120
rect 149 0 195 37
rect 373 83 419 120
rect 373 0 419 37
<< labels >>
flabel metal1 s -52 60 -52 60 0 FreeSans 200 0 0 0 S
flabel metal1 s 396 60 396 60 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 60 172 60 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 421270
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 419800
<< end >>
