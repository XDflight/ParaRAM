magic
tech gf180mcuC
timestamp 1666464484
<< properties >>
string GDS_END 1901258
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1887110
<< end >>
