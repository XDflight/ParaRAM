magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 5014 1094
<< pwell >>
rect -86 -86 5014 453
<< mvnmos >>
rect 124 206 244 324
rect 348 206 468 324
rect 516 206 636 324
rect 740 206 860 324
rect 908 206 1028 324
rect 1362 158 1482 316
rect 1586 158 1706 316
rect 1954 157 2074 275
rect 2178 157 2298 275
rect 2346 157 2466 275
rect 2658 215 2778 333
rect 2862 215 2982 333
rect 3086 215 3206 333
rect 3310 215 3430 333
rect 3826 204 3946 322
rect 3994 204 4114 322
rect 4294 134 4414 292
rect 4662 69 4782 333
<< mvpmos >>
rect 134 644 234 844
rect 348 644 448 844
rect 496 644 596 844
rect 740 644 840 844
rect 900 644 1000 844
rect 1372 577 1472 853
rect 1586 577 1686 853
rect 1964 582 2064 782
rect 2178 582 2278 782
rect 2346 582 2446 782
rect 2658 582 2758 782
rect 2862 582 2962 782
rect 3314 582 3414 782
rect 3518 582 3618 782
rect 3866 592 3966 792
rect 4070 592 4170 792
rect 4314 656 4414 932
rect 4672 574 4772 940
<< mvndiff >>
rect 36 279 124 324
rect 36 233 49 279
rect 95 233 124 279
rect 36 206 124 233
rect 244 279 348 324
rect 244 233 273 279
rect 319 233 348 279
rect 244 206 348 233
rect 468 206 516 324
rect 636 279 740 324
rect 636 233 665 279
rect 711 233 740 279
rect 636 206 740 233
rect 860 206 908 324
rect 1028 206 1150 324
rect 1090 128 1150 206
rect 1274 285 1362 316
rect 1274 239 1287 285
rect 1333 239 1362 285
rect 1274 158 1362 239
rect 1482 217 1586 316
rect 1482 171 1511 217
rect 1557 171 1586 217
rect 1482 158 1586 171
rect 1706 285 1794 316
rect 1706 239 1735 285
rect 1781 239 1794 285
rect 2578 275 2658 333
rect 1706 158 1794 239
rect 1866 216 1954 275
rect 1866 170 1879 216
rect 1925 170 1954 216
rect 1078 115 1150 128
rect 1078 69 1091 115
rect 1137 69 1150 115
rect 1078 56 1150 69
rect 1866 157 1954 170
rect 2074 262 2178 275
rect 2074 216 2103 262
rect 2149 216 2178 262
rect 2074 157 2178 216
rect 2298 157 2346 275
rect 2466 215 2658 275
rect 2778 215 2862 333
rect 2982 320 3086 333
rect 2982 274 3011 320
rect 3057 274 3086 320
rect 2982 215 3086 274
rect 3206 279 3310 333
rect 3206 233 3235 279
rect 3281 233 3310 279
rect 3206 215 3310 233
rect 3430 285 3518 333
rect 3430 239 3459 285
rect 3505 239 3518 285
rect 3430 215 3518 239
rect 2466 157 2598 215
rect 2526 125 2598 157
rect 2526 79 2539 125
rect 2585 79 2598 125
rect 2526 66 2598 79
rect 3738 285 3826 322
rect 3738 239 3751 285
rect 3797 239 3826 285
rect 3738 204 3826 239
rect 3946 204 3994 322
rect 4114 292 4194 322
rect 4114 204 4294 292
rect 4174 134 4294 204
rect 4414 279 4502 292
rect 4414 233 4443 279
rect 4489 233 4502 279
rect 4414 134 4502 233
rect 4574 222 4662 333
rect 4174 124 4234 134
rect 4162 111 4234 124
rect 4162 65 4175 111
rect 4221 65 4234 111
rect 4574 82 4587 222
rect 4633 82 4662 222
rect 4574 69 4662 82
rect 4782 320 4870 333
rect 4782 180 4811 320
rect 4857 180 4870 320
rect 4782 69 4870 180
rect 4162 52 4234 65
<< mvpdiff >>
rect 46 801 134 844
rect 46 661 59 801
rect 105 661 134 801
rect 46 644 134 661
rect 234 831 348 844
rect 234 691 263 831
rect 309 691 348 831
rect 234 644 348 691
rect 448 644 496 844
rect 596 831 740 844
rect 596 691 665 831
rect 711 691 740 831
rect 596 644 740 691
rect 840 644 900 844
rect 1000 801 1088 844
rect 1000 661 1029 801
rect 1075 661 1088 801
rect 1000 644 1088 661
rect 1284 645 1372 853
rect 1284 599 1297 645
rect 1343 599 1372 645
rect 1284 577 1372 599
rect 1472 840 1586 853
rect 1472 794 1501 840
rect 1547 794 1586 840
rect 1472 577 1586 794
rect 1686 636 1774 853
rect 2506 918 2578 931
rect 2506 782 2519 918
rect 1686 590 1715 636
rect 1761 590 1774 636
rect 1686 577 1774 590
rect 1876 737 1964 782
rect 1876 597 1889 737
rect 1935 597 1964 737
rect 1876 582 1964 597
rect 2064 735 2178 782
rect 2064 595 2103 735
rect 2149 595 2178 735
rect 2064 582 2178 595
rect 2278 582 2346 782
rect 2446 778 2519 782
rect 2565 782 2578 918
rect 4226 919 4314 932
rect 4226 873 4239 919
rect 4285 873 4314 919
rect 4226 864 4314 873
rect 4230 792 4314 864
rect 2565 778 2658 782
rect 2446 582 2658 778
rect 2758 641 2862 782
rect 2758 595 2787 641
rect 2833 595 2862 641
rect 2758 582 2862 595
rect 2962 769 3050 782
rect 2962 629 2991 769
rect 3037 629 3050 769
rect 2962 582 3050 629
rect 3226 735 3314 782
rect 3226 595 3239 735
rect 3285 595 3314 735
rect 3226 582 3314 595
rect 3414 769 3518 782
rect 3414 629 3443 769
rect 3489 629 3518 769
rect 3414 582 3518 629
rect 3618 769 3706 782
rect 3618 629 3647 769
rect 3693 629 3706 769
rect 3618 582 3706 629
rect 3778 737 3866 792
rect 3778 691 3791 737
rect 3837 691 3866 737
rect 3778 592 3866 691
rect 3966 779 4070 792
rect 3966 639 3995 779
rect 4041 639 4070 779
rect 3966 592 4070 639
rect 4170 656 4314 792
rect 4414 809 4502 932
rect 4414 669 4443 809
rect 4489 669 4502 809
rect 4414 656 4502 669
rect 4584 801 4672 940
rect 4584 661 4597 801
rect 4643 661 4672 801
rect 4170 592 4250 656
rect 4584 574 4672 661
rect 4772 801 4860 940
rect 4772 661 4801 801
rect 4847 661 4860 801
rect 4772 574 4860 661
<< mvndiffc >>
rect 49 233 95 279
rect 273 233 319 279
rect 665 233 711 279
rect 1287 239 1333 285
rect 1511 171 1557 217
rect 1735 239 1781 285
rect 1879 170 1925 216
rect 1091 69 1137 115
rect 2103 216 2149 262
rect 3011 274 3057 320
rect 3235 233 3281 279
rect 3459 239 3505 285
rect 2539 79 2585 125
rect 3751 239 3797 285
rect 4443 233 4489 279
rect 4175 65 4221 111
rect 4587 82 4633 222
rect 4811 180 4857 320
<< mvpdiffc >>
rect 59 661 105 801
rect 263 691 309 831
rect 665 691 711 831
rect 1029 661 1075 801
rect 1297 599 1343 645
rect 1501 794 1547 840
rect 1715 590 1761 636
rect 1889 597 1935 737
rect 2103 595 2149 735
rect 2519 778 2565 918
rect 4239 873 4285 919
rect 2787 595 2833 641
rect 2991 629 3037 769
rect 3239 595 3285 735
rect 3443 629 3489 769
rect 3647 629 3693 769
rect 3791 691 3837 737
rect 3995 639 4041 779
rect 4443 669 4489 809
rect 4597 661 4643 801
rect 4801 661 4847 801
<< polysilicon >>
rect 134 936 1000 976
rect 134 844 234 936
rect 348 844 448 888
rect 496 844 596 888
rect 740 844 840 888
rect 900 844 1000 936
rect 1586 936 2278 976
rect 1372 853 1472 897
rect 1586 853 1686 936
rect 2178 861 2278 936
rect 134 514 234 644
rect 124 501 234 514
rect 124 455 137 501
rect 183 455 234 501
rect 124 368 234 455
rect 348 501 448 644
rect 348 455 361 501
rect 407 455 448 501
rect 348 368 448 455
rect 496 501 596 644
rect 496 455 509 501
rect 555 455 596 501
rect 496 442 596 455
rect 740 501 840 644
rect 900 600 1000 644
rect 1964 782 2064 826
rect 2178 815 2219 861
rect 2265 815 2278 861
rect 2178 782 2278 815
rect 2346 782 2446 826
rect 2862 922 3966 962
rect 4314 932 4414 976
rect 4672 940 4772 984
rect 2658 782 2758 826
rect 2862 782 2962 922
rect 3314 861 3414 874
rect 3314 815 3327 861
rect 3373 815 3414 861
rect 3314 782 3414 815
rect 3518 782 3618 826
rect 3866 792 3966 922
rect 4070 792 4170 836
rect 1372 514 1472 577
rect 740 455 753 501
rect 799 455 840 501
rect 740 368 840 455
rect 1356 501 1472 514
rect 1356 455 1369 501
rect 1415 455 1472 501
rect 1356 442 1472 455
rect 908 403 1028 416
rect 124 324 244 368
rect 348 324 468 368
rect 516 324 636 368
rect 740 324 860 368
rect 908 357 921 403
rect 967 357 1028 403
rect 908 324 1028 357
rect 1362 360 1472 442
rect 1586 501 1686 577
rect 1586 455 1599 501
rect 1645 455 1686 501
rect 1586 360 1686 455
rect 1964 501 2064 582
rect 2178 538 2278 582
rect 2346 549 2446 582
rect 1964 455 1977 501
rect 2023 490 2064 501
rect 2346 503 2387 549
rect 2433 503 2446 549
rect 2023 455 2298 490
rect 1964 418 2298 455
rect 1362 316 1482 360
rect 1586 316 1706 360
rect 2178 354 2298 418
rect 124 97 244 206
rect 348 162 468 206
rect 516 97 636 206
rect 740 162 860 206
rect 908 162 1028 206
rect 1954 275 2074 319
rect 2178 308 2239 354
rect 2285 308 2298 354
rect 2178 275 2298 308
rect 2346 319 2446 503
rect 2658 457 2758 582
rect 2658 411 2671 457
rect 2717 411 2758 457
rect 2658 377 2758 411
rect 2862 377 2962 582
rect 3314 377 3414 582
rect 3518 538 3618 582
rect 2658 333 2778 377
rect 2862 333 2982 377
rect 3086 333 3206 377
rect 3310 333 3430 377
rect 2346 275 2466 319
rect 124 25 636 97
rect 1362 114 1482 158
rect 1586 97 1706 158
rect 2658 171 2778 215
rect 2862 171 2982 215
rect 3086 182 3206 215
rect 1954 97 2074 157
rect 2178 113 2298 157
rect 2346 113 2466 157
rect 1586 25 2074 97
rect 3086 136 3099 182
rect 3145 136 3206 182
rect 3310 171 3430 215
rect 3086 123 3206 136
rect 3578 123 3618 538
rect 3866 548 3966 592
rect 3866 514 3946 548
rect 3826 501 3946 514
rect 3826 455 3839 501
rect 3885 455 3946 501
rect 3826 322 3946 455
rect 4070 501 4170 592
rect 4070 455 4111 501
rect 4157 455 4170 501
rect 4070 439 4170 455
rect 3994 382 4170 439
rect 4314 501 4414 656
rect 4672 514 4772 574
rect 4314 455 4327 501
rect 4373 455 4414 501
rect 3994 322 4114 382
rect 4314 336 4414 455
rect 4629 501 4772 514
rect 4629 455 4642 501
rect 4688 455 4772 501
rect 4629 442 4772 455
rect 4294 292 4414 336
rect 4662 377 4772 442
rect 4662 333 4782 377
rect 3826 160 3946 204
rect 3994 160 4114 204
rect 3086 51 3618 123
rect 4294 90 4414 134
rect 4662 25 4782 69
<< polycontact >>
rect 137 455 183 501
rect 361 455 407 501
rect 509 455 555 501
rect 2219 815 2265 861
rect 3327 815 3373 861
rect 753 455 799 501
rect 1369 455 1415 501
rect 921 357 967 403
rect 1599 455 1645 501
rect 1977 455 2023 501
rect 2387 503 2433 549
rect 2239 308 2285 354
rect 2671 411 2717 457
rect 3099 136 3145 182
rect 3839 455 3885 501
rect 4111 455 4157 501
rect 4327 455 4373 501
rect 4642 455 4688 501
<< metal1 >>
rect 0 919 4928 1098
rect 0 918 4239 919
rect 263 831 309 918
rect 59 801 105 812
rect 263 680 309 691
rect 665 831 711 842
rect 1029 801 1075 918
rect 711 691 983 726
rect 665 680 983 691
rect 59 634 105 661
rect 59 588 891 634
rect 30 501 194 542
rect 30 455 137 501
rect 183 455 194 501
rect 254 501 418 542
rect 254 455 361 501
rect 407 455 418 501
rect 509 501 555 588
rect 509 409 555 455
rect 49 363 555 409
rect 702 501 799 542
rect 702 455 753 501
rect 49 279 95 363
rect 702 354 799 455
rect 845 414 891 588
rect 937 604 983 680
rect 1490 840 1558 918
rect 1490 794 1501 840
rect 1547 794 1558 840
rect 2219 861 2265 872
rect 1029 650 1075 661
rect 1121 737 1935 748
rect 1121 702 1889 737
rect 1121 604 1167 702
rect 937 558 1167 604
rect 1297 645 1535 656
rect 1343 599 1535 645
rect 1297 588 1535 599
rect 1262 501 1426 542
rect 1262 455 1369 501
rect 1415 455 1426 501
rect 1489 501 1535 588
rect 1715 636 1761 647
rect 1715 501 1761 590
rect 1889 586 1935 597
rect 2103 735 2149 746
rect 2219 721 2265 815
rect 2519 767 2565 778
rect 2991 769 3037 918
rect 2605 721 2945 744
rect 2219 698 2945 721
rect 2219 675 2645 698
rect 1489 455 1599 501
rect 1645 455 1656 501
rect 1715 455 1977 501
rect 2023 455 2034 501
rect 2103 457 2149 595
rect 2787 641 2833 652
rect 2787 549 2833 595
rect 2376 503 2387 549
rect 2433 503 2833 549
rect 2899 572 2945 698
rect 2991 618 3037 629
rect 3147 861 3373 872
rect 3147 815 3327 861
rect 3147 804 3373 815
rect 3147 572 3193 804
rect 3443 769 3489 780
rect 2899 526 3193 572
rect 3239 735 3285 746
rect 845 403 967 414
rect 1489 412 1535 455
rect 1443 409 1535 412
rect 845 357 921 403
rect 845 346 967 357
rect 1287 366 1535 409
rect 1287 363 1460 366
rect 49 222 95 233
rect 273 279 319 290
rect 273 90 319 233
rect 665 279 711 290
rect 665 218 711 233
rect 1287 285 1333 363
rect 1477 317 1649 320
rect 1287 228 1333 239
rect 1379 274 1649 317
rect 1379 271 1494 274
rect 665 182 1242 218
rect 1379 182 1425 271
rect 665 172 1425 182
rect 1197 136 1425 172
rect 1511 217 1557 228
rect 1091 115 1137 126
rect 0 69 1091 90
rect 1511 90 1557 171
rect 1603 182 1649 274
rect 1715 285 1781 455
rect 1715 239 1735 285
rect 1715 228 1781 239
rect 2103 411 2671 457
rect 2717 411 2728 457
rect 2103 262 2149 411
rect 1879 216 1925 227
rect 1603 170 1879 182
rect 2103 205 2149 216
rect 2239 354 2285 365
rect 2239 217 2285 308
rect 2787 309 2833 503
rect 3239 382 3285 595
rect 3443 388 3489 629
rect 3011 336 3285 382
rect 3367 342 3489 388
rect 3634 769 3693 780
rect 3634 629 3647 769
rect 3791 737 3837 918
rect 4285 918 4928 919
rect 4239 862 4285 873
rect 4443 809 4489 820
rect 3791 680 3837 691
rect 3995 779 4041 790
rect 3995 634 4041 639
rect 3693 629 4041 634
rect 3634 588 4041 629
rect 4443 604 4489 669
rect 4597 801 4643 918
rect 4597 650 4643 661
rect 4734 801 4857 812
rect 4734 661 4801 801
rect 4847 661 4857 801
rect 3011 320 3057 336
rect 2787 274 3011 309
rect 2787 263 3057 274
rect 3235 279 3281 290
rect 2239 182 3156 217
rect 2239 171 3099 182
rect 1603 136 1925 170
rect 3088 136 3099 171
rect 3145 136 3156 182
rect 3235 182 3281 233
rect 3367 182 3413 342
rect 3634 296 3680 588
rect 4111 558 4489 604
rect 3726 501 3885 542
rect 3726 455 3839 501
rect 3726 354 3885 455
rect 4111 501 4157 558
rect 4443 512 4489 558
rect 4111 444 4157 455
rect 4327 501 4373 512
rect 3459 285 3797 296
rect 3505 239 3751 285
rect 3459 228 3797 239
rect 4327 214 4373 455
rect 4443 501 4688 512
rect 4443 455 4642 501
rect 4443 444 4688 455
rect 4443 279 4489 444
rect 4734 320 4857 661
rect 4443 222 4489 233
rect 4587 222 4633 233
rect 3841 182 4373 214
rect 3235 168 4373 182
rect 3235 136 3885 168
rect 2528 90 2539 125
rect 1137 79 2539 90
rect 2585 90 2596 125
rect 4175 111 4221 122
rect 2585 79 4175 90
rect 1137 69 4175 79
rect 0 65 4175 69
rect 4221 82 4587 90
rect 4734 180 4811 320
rect 4734 169 4857 180
rect 4633 82 4928 90
rect 4221 65 4928 82
rect 0 -90 4928 65
<< labels >>
flabel metal1 s 1262 455 1426 542 0 FreeSans 200 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 702 354 799 542 0 FreeSans 200 0 0 0 D
port 1 nsew default input
flabel metal1 s 4734 169 4857 812 0 FreeSans 200 0 0 0 Q
port 6 nsew default output
flabel metal1 s 30 455 194 542 0 FreeSans 200 0 0 0 SE
port 2 nsew default input
flabel metal1 s 3726 354 3885 542 0 FreeSans 200 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 254 455 418 542 0 FreeSans 200 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 918 4928 1098 0 FreeSans 200 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 273 233 319 290 0 FreeSans 200 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 4597 862 4643 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4239 862 4285 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3791 862 3837 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 862 3037 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2519 862 2565 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1490 862 1558 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1029 862 1075 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 862 309 918 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4597 794 4643 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3791 794 3837 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 794 3037 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2519 794 2565 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1490 794 1558 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1029 794 1075 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 794 309 862 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4597 767 4643 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3791 767 3837 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 767 3037 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2519 767 2565 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1029 767 1075 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 767 309 794 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4597 680 4643 767 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3791 680 3837 767 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 680 3037 767 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1029 680 1075 767 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 263 680 309 767 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4597 650 4643 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 650 3037 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1029 650 1075 680 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2991 618 3037 650 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4587 228 4633 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 228 319 233 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4587 126 4633 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1511 126 1557 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 126 319 228 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4587 125 4633 126 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1511 125 1557 126 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1091 125 1137 126 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 125 319 126 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4587 122 4633 125 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2528 122 2596 125 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1511 122 1557 125 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1091 122 1137 125 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 122 319 125 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4587 90 4633 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4175 90 4221 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2528 90 2596 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1511 90 1557 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1091 90 1137 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 122 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 4928 90 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4928 1008
string GDS_END 408444
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 397098
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
