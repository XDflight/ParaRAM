magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -58 1371 57 1373
rect -64 1332 64 1371
rect -64 1280 -26 1332
rect 26 1280 64 1332
rect -64 1114 64 1280
rect -64 1062 -26 1114
rect 26 1062 64 1114
rect -64 897 64 1062
rect -64 845 -26 897
rect 26 845 64 897
rect -64 679 64 845
rect -64 627 -26 679
rect 26 627 64 679
rect -64 461 64 627
rect -64 409 -26 461
rect 26 409 64 461
rect -64 244 64 409
rect -64 192 -26 244
rect 26 192 64 244
rect -64 26 64 192
rect -64 -26 -26 26
rect 26 -26 64 26
rect -64 -192 64 -26
rect -64 -244 -26 -192
rect 26 -244 64 -192
rect -64 -409 64 -244
rect -64 -461 -26 -409
rect 26 -461 64 -409
rect -64 -627 64 -461
rect -64 -679 -26 -627
rect 26 -679 64 -627
rect -64 -845 64 -679
rect -64 -897 -26 -845
rect 26 -897 64 -845
rect -64 -1062 64 -897
rect -64 -1091 -26 -1062
rect -65 -1114 -26 -1091
rect 26 -1091 64 -1062
rect 26 -1114 65 -1091
rect -65 -1280 65 -1114
rect -65 -1332 -26 -1280
rect 26 -1332 65 -1280
rect -65 -1373 65 -1332
<< via1 >>
rect -26 1280 26 1332
rect -26 1062 26 1114
rect -26 845 26 897
rect -26 627 26 679
rect -26 409 26 461
rect -26 192 26 244
rect -26 -26 26 26
rect -26 -244 26 -192
rect -26 -461 26 -409
rect -26 -679 26 -627
rect -26 -897 26 -845
rect -26 -1114 26 -1062
rect -26 -1332 26 -1280
<< metal2 >>
rect -64 1332 64 1371
rect -64 1280 -26 1332
rect 26 1280 64 1332
rect -64 1114 64 1280
rect -64 1062 -26 1114
rect 26 1062 64 1114
rect -64 897 64 1062
rect -64 845 -26 897
rect 26 845 64 897
rect -64 679 64 845
rect -64 627 -26 679
rect 26 627 64 679
rect -64 461 64 627
rect -64 409 -26 461
rect 26 409 64 461
rect -64 244 64 409
rect -64 192 -26 244
rect 26 192 64 244
rect -64 26 64 192
rect -64 -26 -26 26
rect 26 -26 64 26
rect -64 -192 64 -26
rect -64 -244 -26 -192
rect 26 -244 64 -192
rect -64 -409 64 -244
rect -64 -461 -26 -409
rect 26 -461 64 -409
rect -64 -627 64 -461
rect -64 -679 -26 -627
rect 26 -679 64 -627
rect -64 -845 64 -679
rect -64 -897 -26 -845
rect 26 -897 64 -845
rect -64 -1062 64 -897
rect -64 -1114 -26 -1062
rect 26 -1114 64 -1062
rect -64 -1280 64 -1114
rect -64 -1332 -26 -1280
rect 26 -1332 64 -1280
rect -64 -1373 64 -1332
<< properties >>
string GDS_END 355062
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 354034
<< end >>
