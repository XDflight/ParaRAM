magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -142 568 894
<< polysilicon >>
rect -31 754 88 826
rect 193 754 312 826
rect -31 -74 88 -1
rect 193 -74 312 -1
use pmos_5p04310589983277_64x8m81  pmos_5p04310589983277_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 552 874
<< properties >>
string GDS_END 753472
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 753030
<< end >>
