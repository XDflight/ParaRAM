magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 29138 51874 56005 52390
rect 29138 50321 32850 51874
rect 35260 50809 39818 51874
rect 35260 50633 39436 50809
rect 45169 50633 49764 51874
rect 52285 50633 56005 51874
<< pwell >>
rect 1774 51482 24710 51514
rect 1774 35138 24710 35170
<< mvpmos >>
rect 7024 32969 7144 33651
rect 7249 32969 7369 33651
rect 7715 32969 7835 33651
rect 7940 32969 8060 33651
rect 17824 32969 17944 33651
rect 18049 32969 18169 33651
rect 18515 32969 18635 33651
rect 18740 32969 18860 33651
rect 66600 32969 66720 33651
rect 66825 32969 66945 33651
rect 67291 32969 67411 33651
rect 67516 32969 67636 33651
rect 77400 32969 77520 33651
rect 77625 32969 77745 33651
rect 78091 32969 78211 33651
rect 78316 32969 78436 33651
rect 7024 32194 7144 32876
rect 7249 32194 7369 32876
rect 7715 32194 7835 32876
rect 7940 32194 8060 32876
rect 17824 32194 17944 32876
rect 18049 32194 18169 32876
rect 18515 32194 18635 32876
rect 18740 32194 18860 32876
rect 66600 32194 66720 32876
rect 66825 32194 66945 32876
rect 67291 32194 67411 32876
rect 67516 32194 67636 32876
rect 77400 32194 77520 32876
rect 77625 32194 77745 32876
rect 78091 32194 78211 32876
rect 78316 32194 78436 32876
<< mvpsubdiff >>
rect 27479 52845 28511 53046
rect 56613 52845 57645 53046
rect 28342 51528 28511 51709
rect 56613 51528 57004 51709
rect 28342 35977 28911 51528
rect 56256 35977 57004 51528
rect 3139 32969 3273 33651
rect 4378 32969 4512 33651
rect 5616 32969 5750 33651
rect 6855 32969 6918 33651
rect 7475 32969 7609 33651
rect 8166 32969 8229 33651
rect 9334 32969 9468 33651
rect 10572 32969 10706 33651
rect 11811 32969 11945 33651
rect 13939 32969 14073 33651
rect 15178 32969 15312 33651
rect 16416 32969 16550 33651
rect 17655 32969 17718 33651
rect 18275 32969 18409 33651
rect 18966 32969 19029 33651
rect 20134 32969 20268 33651
rect 21372 32969 21506 33651
rect 22611 32969 22745 33651
rect 62715 32969 62849 33651
rect 63954 32969 64088 33651
rect 65192 32969 65326 33651
rect 66431 32969 66494 33651
rect 67051 32969 67185 33651
rect 67742 32969 67805 33651
rect 68910 32969 69044 33651
rect 70148 32969 70282 33651
rect 71387 32969 71521 33651
rect 73515 32969 73649 33651
rect 74754 32969 74888 33651
rect 75992 32969 76126 33651
rect 77231 32969 77294 33651
rect 77851 32969 77985 33651
rect 78542 32969 78605 33651
rect 79710 32969 79844 33651
rect 80948 32969 81082 33651
rect 82187 32969 82321 33651
rect 3139 32194 3273 32876
rect 4378 32194 4512 32876
rect 5616 32194 5750 32876
rect 6855 32194 6918 32876
rect 7475 32194 7609 32876
rect 8166 32194 8229 32876
rect 9334 32194 9468 32876
rect 10572 32194 10706 32876
rect 11811 32194 11945 32876
rect 13939 32194 14073 32876
rect 15178 32194 15312 32876
rect 16416 32194 16550 32876
rect 17655 32194 17718 32876
rect 18275 32194 18409 32876
rect 18966 32194 19029 32876
rect 20134 32194 20268 32876
rect 21372 32194 21506 32876
rect 22611 32194 22745 32876
rect 62715 32194 62849 32876
rect 63954 32194 64088 32876
rect 65192 32194 65326 32876
rect 66431 32194 66494 32876
rect 67051 32194 67185 32876
rect 67742 32194 67805 32876
rect 68910 32194 69044 32876
rect 70148 32194 70282 32876
rect 71387 32194 71521 32876
rect 73515 32194 73649 32876
rect 74754 32194 74888 32876
rect 75992 32194 76126 32876
rect 77231 32194 77294 32876
rect 77851 32194 77985 32876
rect 78542 32194 78605 32876
rect 79710 32194 79844 32876
rect 80948 32194 81082 32876
rect 82187 32194 82321 32876
<< metal1 >>
rect 25313 51195 26039 52644
rect 27387 51526 28911 53137
rect 27387 51494 28757 51526
rect 27387 51453 29146 51494
rect 27387 51401 27790 51453
rect 27842 51401 28001 51453
rect 28053 51401 28212 51453
rect 28264 51401 28423 51453
rect 28475 51401 28634 51453
rect 28686 51401 28845 51453
rect 28897 51401 29056 51453
rect 29108 51401 29146 51453
rect 27387 51360 29146 51401
rect 27387 49694 28757 51360
rect 50636 51285 51451 52995
rect 55927 51494 57369 53223
rect 55927 51453 57371 51494
rect 55927 51401 56015 51453
rect 56067 51401 56226 51453
rect 56278 51401 56437 51453
rect 56489 51401 56648 51453
rect 56700 51401 56859 51453
rect 56911 51401 57070 51453
rect 57122 51401 57281 51453
rect 57333 51401 57371 51453
rect 55927 51360 57371 51401
rect 55927 49694 57369 51360
rect 58791 51258 59517 52644
rect 27387 49653 29146 49694
rect 27387 49601 27790 49653
rect 27842 49601 28001 49653
rect 28053 49601 28212 49653
rect 28264 49601 28423 49653
rect 28475 49601 28634 49653
rect 28686 49601 28845 49653
rect 28897 49601 29056 49653
rect 29108 49601 29146 49653
rect 27387 49560 29146 49601
rect 55927 49653 57371 49694
rect 55927 49601 56015 49653
rect 56067 49601 56226 49653
rect 56278 49601 56437 49653
rect 56489 49601 56648 49653
rect 56700 49601 56859 49653
rect 56911 49601 57070 49653
rect 57122 49601 57281 49653
rect 57333 49601 57371 49653
rect 55927 49560 57371 49601
rect 27387 47894 28757 49560
rect 55927 47894 57369 49560
rect 27387 47853 29146 47894
rect 27387 47801 27790 47853
rect 27842 47801 28001 47853
rect 28053 47801 28212 47853
rect 28264 47801 28423 47853
rect 28475 47801 28634 47853
rect 28686 47801 28845 47853
rect 28897 47801 29056 47853
rect 29108 47801 29146 47853
rect 27387 47760 29146 47801
rect 55927 47853 57371 47894
rect 55927 47801 56015 47853
rect 56067 47801 56226 47853
rect 56278 47801 56437 47853
rect 56489 47801 56648 47853
rect 56700 47801 56859 47853
rect 56911 47801 57070 47853
rect 57122 47801 57281 47853
rect 57333 47801 57371 47853
rect 55927 47760 57371 47801
rect 27387 46094 28757 47760
rect 55927 46094 57369 47760
rect 27387 46053 29146 46094
rect 27387 46001 27790 46053
rect 27842 46001 28001 46053
rect 28053 46001 28212 46053
rect 28264 46001 28423 46053
rect 28475 46001 28634 46053
rect 28686 46001 28845 46053
rect 28897 46001 29056 46053
rect 29108 46001 29146 46053
rect 27387 45960 29146 46001
rect 55927 46053 57371 46094
rect 55927 46001 56015 46053
rect 56067 46001 56226 46053
rect 56278 46001 56437 46053
rect 56489 46001 56648 46053
rect 56700 46001 56859 46053
rect 56911 46001 57070 46053
rect 57122 46001 57281 46053
rect 57333 46001 57371 46053
rect 55927 45960 57371 46001
rect 27387 44294 28757 45960
rect 55927 44294 57369 45960
rect 27387 44253 29146 44294
rect 27387 44201 27790 44253
rect 27842 44201 28001 44253
rect 28053 44201 28212 44253
rect 28264 44201 28423 44253
rect 28475 44201 28634 44253
rect 28686 44201 28845 44253
rect 28897 44201 29056 44253
rect 29108 44201 29146 44253
rect 27387 44160 29146 44201
rect 55927 44253 57371 44294
rect 55927 44201 56015 44253
rect 56067 44201 56226 44253
rect 56278 44201 56437 44253
rect 56489 44201 56648 44253
rect 56700 44201 56859 44253
rect 56911 44201 57070 44253
rect 57122 44201 57281 44253
rect 57333 44201 57371 44253
rect 55927 44160 57371 44201
rect 27387 42494 28757 44160
rect 55927 42494 57369 44160
rect 27387 42453 29146 42494
rect 27387 42401 27790 42453
rect 27842 42401 28001 42453
rect 28053 42401 28212 42453
rect 28264 42401 28423 42453
rect 28475 42401 28634 42453
rect 28686 42401 28845 42453
rect 28897 42401 29056 42453
rect 29108 42401 29146 42453
rect 27387 42360 29146 42401
rect 55927 42453 57371 42494
rect 55927 42401 56015 42453
rect 56067 42401 56226 42453
rect 56278 42401 56437 42453
rect 56489 42401 56648 42453
rect 56700 42401 56859 42453
rect 56911 42401 57070 42453
rect 57122 42401 57281 42453
rect 57333 42401 57371 42453
rect 55927 42360 57371 42401
rect 27387 40694 28757 42360
rect 55927 40694 57369 42360
rect 27387 40653 29146 40694
rect 27387 40601 27790 40653
rect 27842 40601 28001 40653
rect 28053 40601 28212 40653
rect 28264 40601 28423 40653
rect 28475 40601 28634 40653
rect 28686 40601 28845 40653
rect 28897 40601 29056 40653
rect 29108 40601 29146 40653
rect 27387 40560 29146 40601
rect 55927 40653 57371 40694
rect 55927 40601 56015 40653
rect 56067 40601 56226 40653
rect 56278 40601 56437 40653
rect 56489 40601 56648 40653
rect 56700 40601 56859 40653
rect 56911 40601 57070 40653
rect 57122 40601 57281 40653
rect 57333 40601 57371 40653
rect 55927 40560 57371 40601
rect 27387 38894 28757 40560
rect 55927 38894 57369 40560
rect 27387 38853 29146 38894
rect 27387 38801 27790 38853
rect 27842 38801 28001 38853
rect 28053 38801 28212 38853
rect 28264 38801 28423 38853
rect 28475 38801 28634 38853
rect 28686 38801 28845 38853
rect 28897 38801 29056 38853
rect 29108 38801 29146 38853
rect 27387 38760 29146 38801
rect 55927 38853 57371 38894
rect 55927 38801 56015 38853
rect 56067 38801 56226 38853
rect 56278 38801 56437 38853
rect 56489 38801 56648 38853
rect 56700 38801 56859 38853
rect 56911 38801 57070 38853
rect 57122 38801 57281 38853
rect 57333 38801 57371 38853
rect 55927 38760 57371 38801
rect 27387 37094 28757 38760
rect 55927 37094 57369 38760
rect 27387 37053 29146 37094
rect 27387 37001 27790 37053
rect 27842 37001 28001 37053
rect 28053 37001 28212 37053
rect 28264 37001 28423 37053
rect 28475 37001 28634 37053
rect 28686 37001 28845 37053
rect 28897 37001 29056 37053
rect 29108 37001 29146 37053
rect 27387 36960 29146 37001
rect 55927 37053 57371 37094
rect 55927 37001 56015 37053
rect 56067 37001 56226 37053
rect 56278 37001 56437 37053
rect 56489 37001 56648 37053
rect 56700 37001 56859 37053
rect 56911 37001 57070 37053
rect 57122 37001 57281 37053
rect 57333 37001 57371 37053
rect 55927 36960 57371 37001
rect 27387 35985 28757 36960
rect 55927 35985 57369 36960
rect 27387 34613 27828 35985
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 84369 35126 85931 35326
rect 27387 34245 57297 34613
rect 85090 34536 85931 35126
rect 26772 1777 27214 33519
rect 2562 1689 2742 1701
rect 2562 1637 2574 1689
rect 2730 1637 2742 1689
rect 2562 1625 2742 1637
rect 12627 1689 12807 1701
rect 12627 1637 12639 1689
rect 12795 1637 12807 1689
rect 12627 1625 12807 1637
rect 13077 1689 13257 1701
rect 13077 1637 13089 1689
rect 13245 1637 13257 1689
rect 13077 1625 13257 1637
rect 23427 1689 23607 1701
rect 23427 1637 23439 1689
rect 23595 1637 23607 1689
rect 23427 1625 23607 1637
rect 27387 1282 27828 34245
rect 49896 6349 50076 6361
rect 49896 6347 49908 6349
rect 49728 6301 49908 6347
rect 49896 6297 49908 6301
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 57295 5220 57736 33519
rect 57909 5220 58351 33519
rect 83398 32048 83834 32122
rect 51642 5199 51822 5211
rect 51642 5196 51654 5199
rect 49963 5150 51654 5196
rect 51642 5147 51654 5150
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 40610 4904 40790 4916
rect 40610 4852 40622 4904
rect 40778 4852 40790 4904
rect 40610 4840 40790 4852
rect 57295 3584 57736 4728
rect 28628 1282 40180 1666
rect 50834 1282 56586 1662
rect 57295 1282 57737 3584
rect 57909 1777 58351 4728
rect 62138 1689 62318 1701
rect 62138 1637 62150 1689
rect 62306 1637 62318 1689
rect 62138 1625 62318 1637
rect 72203 1689 72383 1701
rect 72203 1637 72215 1689
rect 72371 1637 72383 1689
rect 72203 1625 72383 1637
rect 72653 1689 72833 1701
rect 72653 1637 72665 1689
rect 72821 1637 72833 1689
rect 72653 1625 72833 1637
rect 82718 1689 82898 1701
rect 82718 1637 82730 1689
rect 82886 1637 82898 1689
rect 82718 1625 82898 1637
rect 282 915 86090 1282
rect 282 655 29090 915
rect 29142 655 29792 915
rect 29844 655 86090 915
rect 282 282 86090 655
<< via1 >>
rect 27790 51401 27842 51453
rect 28001 51401 28053 51453
rect 28212 51401 28264 51453
rect 28423 51401 28475 51453
rect 28634 51401 28686 51453
rect 28845 51401 28897 51453
rect 29056 51401 29108 51453
rect 56015 51401 56067 51453
rect 56226 51401 56278 51453
rect 56437 51401 56489 51453
rect 56648 51401 56700 51453
rect 56859 51401 56911 51453
rect 57070 51401 57122 51453
rect 57281 51401 57333 51453
rect 27790 49601 27842 49653
rect 28001 49601 28053 49653
rect 28212 49601 28264 49653
rect 28423 49601 28475 49653
rect 28634 49601 28686 49653
rect 28845 49601 28897 49653
rect 29056 49601 29108 49653
rect 56015 49601 56067 49653
rect 56226 49601 56278 49653
rect 56437 49601 56489 49653
rect 56648 49601 56700 49653
rect 56859 49601 56911 49653
rect 57070 49601 57122 49653
rect 57281 49601 57333 49653
rect 27790 47801 27842 47853
rect 28001 47801 28053 47853
rect 28212 47801 28264 47853
rect 28423 47801 28475 47853
rect 28634 47801 28686 47853
rect 28845 47801 28897 47853
rect 29056 47801 29108 47853
rect 56015 47801 56067 47853
rect 56226 47801 56278 47853
rect 56437 47801 56489 47853
rect 56648 47801 56700 47853
rect 56859 47801 56911 47853
rect 57070 47801 57122 47853
rect 57281 47801 57333 47853
rect 27790 46001 27842 46053
rect 28001 46001 28053 46053
rect 28212 46001 28264 46053
rect 28423 46001 28475 46053
rect 28634 46001 28686 46053
rect 28845 46001 28897 46053
rect 29056 46001 29108 46053
rect 56015 46001 56067 46053
rect 56226 46001 56278 46053
rect 56437 46001 56489 46053
rect 56648 46001 56700 46053
rect 56859 46001 56911 46053
rect 57070 46001 57122 46053
rect 57281 46001 57333 46053
rect 27790 44201 27842 44253
rect 28001 44201 28053 44253
rect 28212 44201 28264 44253
rect 28423 44201 28475 44253
rect 28634 44201 28686 44253
rect 28845 44201 28897 44253
rect 29056 44201 29108 44253
rect 56015 44201 56067 44253
rect 56226 44201 56278 44253
rect 56437 44201 56489 44253
rect 56648 44201 56700 44253
rect 56859 44201 56911 44253
rect 57070 44201 57122 44253
rect 57281 44201 57333 44253
rect 27790 42401 27842 42453
rect 28001 42401 28053 42453
rect 28212 42401 28264 42453
rect 28423 42401 28475 42453
rect 28634 42401 28686 42453
rect 28845 42401 28897 42453
rect 29056 42401 29108 42453
rect 56015 42401 56067 42453
rect 56226 42401 56278 42453
rect 56437 42401 56489 42453
rect 56648 42401 56700 42453
rect 56859 42401 56911 42453
rect 57070 42401 57122 42453
rect 57281 42401 57333 42453
rect 27790 40601 27842 40653
rect 28001 40601 28053 40653
rect 28212 40601 28264 40653
rect 28423 40601 28475 40653
rect 28634 40601 28686 40653
rect 28845 40601 28897 40653
rect 29056 40601 29108 40653
rect 56015 40601 56067 40653
rect 56226 40601 56278 40653
rect 56437 40601 56489 40653
rect 56648 40601 56700 40653
rect 56859 40601 56911 40653
rect 57070 40601 57122 40653
rect 57281 40601 57333 40653
rect 27790 38801 27842 38853
rect 28001 38801 28053 38853
rect 28212 38801 28264 38853
rect 28423 38801 28475 38853
rect 28634 38801 28686 38853
rect 28845 38801 28897 38853
rect 29056 38801 29108 38853
rect 56015 38801 56067 38853
rect 56226 38801 56278 38853
rect 56437 38801 56489 38853
rect 56648 38801 56700 38853
rect 56859 38801 56911 38853
rect 57070 38801 57122 38853
rect 57281 38801 57333 38853
rect 27790 37001 27842 37053
rect 28001 37001 28053 37053
rect 28212 37001 28264 37053
rect 28423 37001 28475 37053
rect 28634 37001 28686 37053
rect 28845 37001 28897 37053
rect 29056 37001 29108 37053
rect 56015 37001 56067 37053
rect 56226 37001 56278 37053
rect 56437 37001 56489 37053
rect 56648 37001 56700 37053
rect 56859 37001 56911 37053
rect 57070 37001 57122 37053
rect 57281 37001 57333 37053
rect 60575 35338 60627 35494
rect 2574 1637 2730 1689
rect 12639 1637 12795 1689
rect 13089 1637 13245 1689
rect 23439 1637 23595 1689
rect 49908 6297 50064 6349
rect 51654 5147 51810 5199
rect 40622 4852 40778 4904
rect 62150 1637 62306 1689
rect 72215 1637 72371 1689
rect 72665 1637 72821 1689
rect 82730 1637 82886 1689
rect 29090 655 29142 915
rect 29792 655 29844 915
<< metal2 >>
rect 282 53168 86090 53494
rect 706 51976 85666 52976
rect 25313 26433 26039 51627
rect 26823 32088 27163 51976
rect 26823 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 27163 32088
rect 26823 31870 27163 32032
rect 26823 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 27163 31870
rect 26823 31652 27163 31814
rect 26823 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 27163 31652
rect 26823 27382 27163 31596
rect 27387 51455 29146 51494
rect 27387 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 29146 51455
rect 27387 51360 29146 51399
rect 27387 49694 27828 51360
rect 29486 51285 30364 51976
rect 30769 51285 32888 51976
rect 35128 51285 36415 51976
rect 38953 51471 39618 51976
rect 48789 51285 49990 51976
rect 52226 51285 54354 51976
rect 54758 51285 55638 51976
rect 55977 51455 57371 51494
rect 55977 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 57371 51455
rect 55977 51360 57371 51399
rect 41865 50613 42045 50623
rect 41865 50453 41875 50613
rect 42035 50453 42045 50613
rect 41865 50443 42045 50453
rect 27387 49655 29146 49694
rect 27387 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 29146 49655
rect 27387 49560 29146 49599
rect 55977 49655 57371 49694
rect 55977 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 57371 49655
rect 55977 49560 57371 49599
rect 27387 47894 27828 49560
rect 27387 47855 29146 47894
rect 27387 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 29146 47855
rect 27387 47760 29146 47799
rect 55977 47855 57371 47894
rect 55977 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 57371 47855
rect 55977 47760 57371 47799
rect 27387 46094 27828 47760
rect 27387 46055 29146 46094
rect 27387 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 29146 46055
rect 27387 45960 29146 45999
rect 55977 46055 57371 46094
rect 55977 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 57371 46055
rect 55977 45960 57371 45999
rect 27387 44294 27828 45960
rect 27387 44255 29146 44294
rect 27387 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 29146 44255
rect 27387 44160 29146 44199
rect 55977 44255 57371 44294
rect 55977 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 57371 44255
rect 55977 44160 57371 44199
rect 27387 42494 27828 44160
rect 27387 42455 29146 42494
rect 27387 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 29146 42455
rect 27387 42360 29146 42399
rect 55977 42455 57371 42494
rect 55977 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 57371 42455
rect 55977 42360 57371 42399
rect 27387 40694 27828 42360
rect 27387 40655 29146 40694
rect 27387 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 29146 40655
rect 27387 40560 29146 40599
rect 55977 40655 57371 40694
rect 55977 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 57371 40655
rect 55977 40560 57371 40599
rect 27387 38894 27828 40560
rect 27387 38855 29146 38894
rect 27387 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 29146 38855
rect 27387 38760 29146 38799
rect 55977 38855 57371 38894
rect 55977 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 57371 38855
rect 55977 38760 57371 38799
rect 27387 37094 27828 38760
rect 27387 37055 29146 37094
rect 27387 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 29146 37055
rect 27387 36960 29146 36999
rect 55977 37055 57371 37094
rect 55977 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 57371 37055
rect 55977 36960 57371 36999
rect 27387 26799 27828 36960
rect 36863 35881 37743 36650
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 36863 35786 37743 35825
rect 41472 35761 41694 36096
rect 38596 35532 41694 35761
rect 38596 35516 38817 35532
rect 31615 35287 38817 35516
rect 41850 35425 42072 35528
rect 31615 33349 31836 35287
rect 39077 35197 42072 35425
rect 39077 35171 39298 35197
rect 31970 34943 39298 35171
rect 42228 35090 42449 36096
rect 31970 33349 32192 34943
rect 39755 34861 42449 35090
rect 39755 34675 39977 34861
rect 42603 34754 42825 36085
rect 38301 34491 39977 34675
rect 37201 34446 39977 34491
rect 40106 34526 42825 34754
rect 37201 34263 38523 34446
rect 40106 34312 40328 34526
rect 42983 34419 43205 36096
rect 37201 33360 37423 34263
rect 38642 34156 40328 34312
rect 37557 34084 40328 34156
rect 40458 34190 43205 34419
rect 37557 33927 38863 34084
rect 40458 33977 40679 34190
rect 43359 34083 43580 36085
rect 45513 35842 45735 36096
rect 37557 33349 37778 33927
rect 38993 33748 40679 33977
rect 40809 33855 43580 34083
rect 44646 35614 45735 35842
rect 38993 33360 39215 33748
rect 40809 33625 41031 33855
rect 39349 33397 41031 33625
rect 44646 33576 44867 35614
rect 45891 35507 46112 36096
rect 44997 35278 46112 35507
rect 46268 35681 46490 36096
rect 46268 35453 46501 35681
rect 44997 33576 45219 35278
rect 46279 33576 46501 35453
rect 46646 35346 46868 36085
rect 46631 35117 46868 35346
rect 46631 33564 46852 35117
rect 47026 34836 47248 36085
rect 47402 35171 47623 36096
rect 47779 35507 48001 36096
rect 48157 35842 48379 36096
rect 48157 35614 50120 35842
rect 47779 35278 49769 35507
rect 47402 34943 48486 35171
rect 47026 34607 48135 34836
rect 47913 33564 48135 34607
rect 48265 33576 48486 34943
rect 49547 33576 49769 35278
rect 49898 33576 50120 35614
rect 27387 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 27387 26581 27828 26743
rect 27387 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 26435 26286 26643 26321
rect 26435 26126 26450 26286
rect 26610 26126 26643 26286
rect 26077 25967 26285 26002
rect 26077 25807 26092 25967
rect 26252 25807 26285 25967
rect 25741 25647 25949 25676
rect 25741 25487 25756 25647
rect 25916 25487 25949 25647
rect 25406 25328 25614 25357
rect 25406 25168 25421 25328
rect 25581 25168 25614 25328
rect 25066 24637 25274 24666
rect 25066 24477 25081 24637
rect 25241 24477 25274 24637
rect 24729 24316 24937 24345
rect 24729 24156 24744 24316
rect 24904 24156 24937 24316
rect 24401 23995 24609 24024
rect 24401 23835 24416 23995
rect 24576 23835 24609 23995
rect 24042 23673 24250 23702
rect 24042 23513 24057 23673
rect 24217 23513 24250 23673
rect 24042 17317 24250 23513
rect 24401 17656 24609 23835
rect 24729 17977 24937 24156
rect 25066 18350 25274 24477
rect 25406 18684 25614 25168
rect 25741 19027 25949 25487
rect 26077 19347 26285 25807
rect 26435 19692 26643 26126
rect 27387 25028 27828 26525
rect 27387 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 27828 25028
rect 27387 24810 27828 24972
rect 27387 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 27828 24810
rect 26914 20570 27094 20580
rect 26914 20410 26924 20570
rect 27084 20410 27094 20570
rect 26914 20400 27094 20410
rect 26914 20226 27094 20236
rect 26914 20066 26924 20226
rect 27084 20066 27094 20226
rect 26914 20056 27094 20066
rect 26435 19532 26465 19692
rect 26625 19532 26643 19692
rect 26435 19502 26643 19532
rect 26077 19187 26107 19347
rect 26267 19187 26285 19347
rect 26077 19162 26285 19187
rect 25741 18867 25771 19027
rect 25931 18867 25949 19027
rect 25741 18822 25949 18867
rect 25406 18524 25434 18684
rect 25594 18524 25614 18684
rect 25406 18482 25614 18524
rect 25066 18190 25094 18350
rect 25254 18190 25274 18350
rect 25066 18142 25274 18190
rect 24729 17817 24757 17977
rect 24917 17817 24937 17977
rect 24729 17803 24937 17817
rect 24401 17496 24429 17656
rect 24589 17496 24609 17656
rect 24401 17462 24609 17496
rect 24042 17157 24069 17317
rect 24229 17157 24250 17317
rect 24042 17122 24250 17157
rect 27387 7535 27828 24754
rect 57295 26799 57736 33519
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 57736 26799
rect 57295 26581 57736 26743
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 57736 26581
rect 51756 9971 51832 9981
rect 51756 9811 51766 9971
rect 51822 9811 51832 9971
rect 51756 9801 51832 9811
rect 49896 8956 50076 8966
rect 49896 8900 49906 8956
rect 50066 8900 50076 8956
rect 49896 8890 50076 8900
rect 27387 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 27387 7317 27828 7479
rect 27387 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 27387 7099 27828 7261
rect 27387 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 27387 6120 27828 7043
rect 49958 6361 50014 8890
rect 49896 6349 50076 6361
rect 49896 6297 49908 6349
rect 50064 6297 50076 6349
rect 49896 6285 50076 6297
rect 27387 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 27828 6120
rect 27387 5902 27828 6064
rect 27387 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 27828 5902
rect 26823 5539 27163 5578
rect 26823 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27163 5539
rect 26823 5321 27163 5483
rect 26823 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27163 5321
rect 26823 5226 27163 5265
rect 1864 5024 2509 5135
rect 11727 5073 11783 5140
rect 1864 0 2088 5024
rect 3263 5001 3357 5062
rect 11617 5017 11783 5073
rect 3263 4880 3604 5001
rect 2539 1689 2763 1701
rect 2539 1637 2574 1689
rect 2730 1637 2763 1689
rect 2539 0 2763 1637
rect 3380 0 3604 4880
rect 11617 1701 11673 5017
rect 12575 4740 12631 5185
rect 12290 4684 12631 4740
rect 13253 4740 13309 5185
rect 14101 5073 14157 5140
rect 14101 5017 14267 5073
rect 13253 4684 13594 4740
rect 12290 1701 12346 4684
rect 13538 1701 13594 4684
rect 14211 1701 14267 5017
rect 22527 5001 22621 5062
rect 23375 5024 24019 5135
rect 22279 4880 22621 5001
rect 11533 0 11757 1701
rect 12206 0 12430 1701
rect 12604 1689 12828 1701
rect 12604 1637 12639 1689
rect 12795 1637 12828 1689
rect 12604 0 12828 1637
rect 13054 1689 13278 1701
rect 13054 1637 13089 1689
rect 13245 1637 13278 1689
rect 13054 0 13278 1637
rect 13454 0 13678 1701
rect 14127 0 14351 1701
rect 22279 0 22503 4880
rect 23404 1689 23628 1701
rect 23404 1637 23439 1689
rect 23595 1637 23628 1689
rect 23404 0 23628 1637
rect 23795 0 24019 5024
rect 26823 4528 27163 4567
rect 26823 4472 26859 4528
rect 26915 4472 27071 4528
rect 27127 4472 27163 4528
rect 26823 4310 27163 4472
rect 26823 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 27163 4310
rect 26823 4215 27163 4254
rect 27387 3837 27828 5846
rect 51766 5211 51822 9801
rect 51642 5199 51822 5211
rect 51642 5147 51654 5199
rect 51810 5147 51822 5199
rect 51642 5135 51822 5147
rect 57295 6120 57736 26525
rect 57295 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 57736 6120
rect 57295 5902 57736 6064
rect 57295 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 57736 5902
rect 40588 4904 40812 4928
rect 40588 4852 40622 4904
rect 40778 4852 40812 4904
rect 27387 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 27828 3837
rect 27387 3619 27828 3781
rect 27387 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 27828 3619
rect 27387 3524 27828 3563
rect 28764 3837 28894 3876
rect 28764 3781 28801 3837
rect 28857 3781 28894 3837
rect 28764 3619 28894 3781
rect 28764 3563 28801 3619
rect 28857 3563 28894 3619
rect 28764 3525 28894 3563
rect 27936 0 28160 3418
rect 29006 3050 29135 3418
rect 29247 3231 29929 3418
rect 29006 915 29230 3050
rect 29006 655 29090 915
rect 29142 655 29230 915
rect 29006 0 29230 655
rect 29705 915 29929 3231
rect 29705 655 29792 915
rect 29844 655 29929 915
rect 29705 0 29929 655
rect 30859 0 31083 3605
rect 32552 0 32776 3605
rect 34243 0 34467 3605
rect 40588 0 40812 4852
rect 43790 3044 43970 3054
rect 43790 2988 43800 3044
rect 43960 2988 43970 3044
rect 43790 2978 43970 2988
rect 48644 282 48997 3873
rect 49145 1232 49498 4618
rect 57295 3837 57736 5846
rect 57295 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 57736 3837
rect 57295 3619 57736 3781
rect 57295 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 57736 3619
rect 57295 3524 57736 3563
rect 57909 32088 58351 51976
rect 57909 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 57909 31870 58351 32032
rect 57909 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 57909 31652 58351 31814
rect 57909 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 57909 20570 58351 31596
rect 58791 26433 59517 51591
rect 60563 35494 60639 35506
rect 60563 35338 60575 35494
rect 60627 35338 60639 35494
rect 60563 35326 60639 35338
rect 57909 20410 58048 20570
rect 58208 20410 58351 20570
rect 57909 20226 58351 20410
rect 57909 20066 58048 20226
rect 58208 20066 58351 20226
rect 57909 5539 58351 20066
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 58351 5539
rect 57909 5321 58351 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 58351 5321
rect 57909 4528 58351 5265
rect 57909 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4472 58351 4528
rect 57909 4310 58351 4472
rect 57909 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 58351 4310
rect 57909 3524 58351 4254
rect 61507 5024 62085 5135
rect 71303 5073 71359 5140
rect 50342 0 50566 3517
rect 53772 3255 55669 3418
rect 53772 0 53996 3255
rect 55781 2974 55911 3418
rect 54417 2789 55911 2974
rect 54417 0 54641 2789
rect 56023 2480 56152 3418
rect 55164 2224 56152 2480
rect 55164 0 55388 2224
rect 56265 0 56489 3481
rect 61507 1701 61601 5024
rect 62839 5001 62933 5062
rect 71193 5017 71359 5073
rect 62839 4880 63115 5001
rect 63021 1701 63115 4880
rect 71193 1701 71249 5017
rect 72151 4740 72207 5185
rect 71866 4684 72207 4740
rect 72829 4740 72885 5185
rect 73677 5073 73733 5140
rect 73677 5017 73843 5073
rect 72829 4684 73170 4740
rect 71866 1701 71922 4684
rect 73114 1701 73170 4684
rect 73787 1701 73843 5017
rect 82103 5001 82197 5062
rect 82951 5024 83529 5135
rect 81921 4880 82197 5001
rect 81921 1701 82015 4880
rect 83435 1701 83529 5024
rect 61447 0 61671 1701
rect 62115 1689 62339 1701
rect 62115 1637 62150 1689
rect 62306 1637 62339 1689
rect 62115 0 62339 1637
rect 62958 0 63182 1701
rect 71109 0 71333 1701
rect 71782 0 72006 1701
rect 72180 1689 72404 1701
rect 72180 1637 72215 1689
rect 72371 1637 72404 1689
rect 72180 0 72404 1637
rect 72630 1689 72854 1701
rect 72630 1637 72665 1689
rect 72821 1637 72854 1689
rect 72630 0 72854 1637
rect 73030 0 73254 1701
rect 73703 0 73927 1701
rect 81855 0 82079 1701
rect 82695 1689 82919 1701
rect 82695 1637 82730 1689
rect 82886 1637 82919 1689
rect 82695 0 82919 1637
rect 83372 0 83596 1701
<< via2 >>
rect 26859 32032 26915 32088
rect 27071 32032 27127 32088
rect 26859 31814 26915 31870
rect 27071 31814 27127 31870
rect 26859 31596 26915 31652
rect 27071 31596 27127 31652
rect 27788 51453 27844 51455
rect 27788 51401 27790 51453
rect 27790 51401 27842 51453
rect 27842 51401 27844 51453
rect 27788 51399 27844 51401
rect 27999 51453 28055 51455
rect 27999 51401 28001 51453
rect 28001 51401 28053 51453
rect 28053 51401 28055 51453
rect 27999 51399 28055 51401
rect 28210 51453 28266 51455
rect 28210 51401 28212 51453
rect 28212 51401 28264 51453
rect 28264 51401 28266 51453
rect 28210 51399 28266 51401
rect 28421 51453 28477 51455
rect 28421 51401 28423 51453
rect 28423 51401 28475 51453
rect 28475 51401 28477 51453
rect 28421 51399 28477 51401
rect 28632 51453 28688 51455
rect 28632 51401 28634 51453
rect 28634 51401 28686 51453
rect 28686 51401 28688 51453
rect 28632 51399 28688 51401
rect 28843 51453 28899 51455
rect 28843 51401 28845 51453
rect 28845 51401 28897 51453
rect 28897 51401 28899 51453
rect 28843 51399 28899 51401
rect 29054 51453 29110 51455
rect 29054 51401 29056 51453
rect 29056 51401 29108 51453
rect 29108 51401 29110 51453
rect 29054 51399 29110 51401
rect 56013 51453 56069 51455
rect 56013 51401 56015 51453
rect 56015 51401 56067 51453
rect 56067 51401 56069 51453
rect 56013 51399 56069 51401
rect 56224 51453 56280 51455
rect 56224 51401 56226 51453
rect 56226 51401 56278 51453
rect 56278 51401 56280 51453
rect 56224 51399 56280 51401
rect 56435 51453 56491 51455
rect 56435 51401 56437 51453
rect 56437 51401 56489 51453
rect 56489 51401 56491 51453
rect 56435 51399 56491 51401
rect 56646 51453 56702 51455
rect 56646 51401 56648 51453
rect 56648 51401 56700 51453
rect 56700 51401 56702 51453
rect 56646 51399 56702 51401
rect 56857 51453 56913 51455
rect 56857 51401 56859 51453
rect 56859 51401 56911 51453
rect 56911 51401 56913 51453
rect 56857 51399 56913 51401
rect 57068 51453 57124 51455
rect 57068 51401 57070 51453
rect 57070 51401 57122 51453
rect 57122 51401 57124 51453
rect 57068 51399 57124 51401
rect 57279 51453 57335 51455
rect 57279 51401 57281 51453
rect 57281 51401 57333 51453
rect 57333 51401 57335 51453
rect 57279 51399 57335 51401
rect 41875 50453 42035 50613
rect 27788 49653 27844 49655
rect 27788 49601 27790 49653
rect 27790 49601 27842 49653
rect 27842 49601 27844 49653
rect 27788 49599 27844 49601
rect 27999 49653 28055 49655
rect 27999 49601 28001 49653
rect 28001 49601 28053 49653
rect 28053 49601 28055 49653
rect 27999 49599 28055 49601
rect 28210 49653 28266 49655
rect 28210 49601 28212 49653
rect 28212 49601 28264 49653
rect 28264 49601 28266 49653
rect 28210 49599 28266 49601
rect 28421 49653 28477 49655
rect 28421 49601 28423 49653
rect 28423 49601 28475 49653
rect 28475 49601 28477 49653
rect 28421 49599 28477 49601
rect 28632 49653 28688 49655
rect 28632 49601 28634 49653
rect 28634 49601 28686 49653
rect 28686 49601 28688 49653
rect 28632 49599 28688 49601
rect 28843 49653 28899 49655
rect 28843 49601 28845 49653
rect 28845 49601 28897 49653
rect 28897 49601 28899 49653
rect 28843 49599 28899 49601
rect 29054 49653 29110 49655
rect 29054 49601 29056 49653
rect 29056 49601 29108 49653
rect 29108 49601 29110 49653
rect 29054 49599 29110 49601
rect 56013 49653 56069 49655
rect 56013 49601 56015 49653
rect 56015 49601 56067 49653
rect 56067 49601 56069 49653
rect 56013 49599 56069 49601
rect 56224 49653 56280 49655
rect 56224 49601 56226 49653
rect 56226 49601 56278 49653
rect 56278 49601 56280 49653
rect 56224 49599 56280 49601
rect 56435 49653 56491 49655
rect 56435 49601 56437 49653
rect 56437 49601 56489 49653
rect 56489 49601 56491 49653
rect 56435 49599 56491 49601
rect 56646 49653 56702 49655
rect 56646 49601 56648 49653
rect 56648 49601 56700 49653
rect 56700 49601 56702 49653
rect 56646 49599 56702 49601
rect 56857 49653 56913 49655
rect 56857 49601 56859 49653
rect 56859 49601 56911 49653
rect 56911 49601 56913 49653
rect 56857 49599 56913 49601
rect 57068 49653 57124 49655
rect 57068 49601 57070 49653
rect 57070 49601 57122 49653
rect 57122 49601 57124 49653
rect 57068 49599 57124 49601
rect 57279 49653 57335 49655
rect 57279 49601 57281 49653
rect 57281 49601 57333 49653
rect 57333 49601 57335 49653
rect 57279 49599 57335 49601
rect 27788 47853 27844 47855
rect 27788 47801 27790 47853
rect 27790 47801 27842 47853
rect 27842 47801 27844 47853
rect 27788 47799 27844 47801
rect 27999 47853 28055 47855
rect 27999 47801 28001 47853
rect 28001 47801 28053 47853
rect 28053 47801 28055 47853
rect 27999 47799 28055 47801
rect 28210 47853 28266 47855
rect 28210 47801 28212 47853
rect 28212 47801 28264 47853
rect 28264 47801 28266 47853
rect 28210 47799 28266 47801
rect 28421 47853 28477 47855
rect 28421 47801 28423 47853
rect 28423 47801 28475 47853
rect 28475 47801 28477 47853
rect 28421 47799 28477 47801
rect 28632 47853 28688 47855
rect 28632 47801 28634 47853
rect 28634 47801 28686 47853
rect 28686 47801 28688 47853
rect 28632 47799 28688 47801
rect 28843 47853 28899 47855
rect 28843 47801 28845 47853
rect 28845 47801 28897 47853
rect 28897 47801 28899 47853
rect 28843 47799 28899 47801
rect 29054 47853 29110 47855
rect 29054 47801 29056 47853
rect 29056 47801 29108 47853
rect 29108 47801 29110 47853
rect 29054 47799 29110 47801
rect 56013 47853 56069 47855
rect 56013 47801 56015 47853
rect 56015 47801 56067 47853
rect 56067 47801 56069 47853
rect 56013 47799 56069 47801
rect 56224 47853 56280 47855
rect 56224 47801 56226 47853
rect 56226 47801 56278 47853
rect 56278 47801 56280 47853
rect 56224 47799 56280 47801
rect 56435 47853 56491 47855
rect 56435 47801 56437 47853
rect 56437 47801 56489 47853
rect 56489 47801 56491 47853
rect 56435 47799 56491 47801
rect 56646 47853 56702 47855
rect 56646 47801 56648 47853
rect 56648 47801 56700 47853
rect 56700 47801 56702 47853
rect 56646 47799 56702 47801
rect 56857 47853 56913 47855
rect 56857 47801 56859 47853
rect 56859 47801 56911 47853
rect 56911 47801 56913 47853
rect 56857 47799 56913 47801
rect 57068 47853 57124 47855
rect 57068 47801 57070 47853
rect 57070 47801 57122 47853
rect 57122 47801 57124 47853
rect 57068 47799 57124 47801
rect 57279 47853 57335 47855
rect 57279 47801 57281 47853
rect 57281 47801 57333 47853
rect 57333 47801 57335 47853
rect 57279 47799 57335 47801
rect 27788 46053 27844 46055
rect 27788 46001 27790 46053
rect 27790 46001 27842 46053
rect 27842 46001 27844 46053
rect 27788 45999 27844 46001
rect 27999 46053 28055 46055
rect 27999 46001 28001 46053
rect 28001 46001 28053 46053
rect 28053 46001 28055 46053
rect 27999 45999 28055 46001
rect 28210 46053 28266 46055
rect 28210 46001 28212 46053
rect 28212 46001 28264 46053
rect 28264 46001 28266 46053
rect 28210 45999 28266 46001
rect 28421 46053 28477 46055
rect 28421 46001 28423 46053
rect 28423 46001 28475 46053
rect 28475 46001 28477 46053
rect 28421 45999 28477 46001
rect 28632 46053 28688 46055
rect 28632 46001 28634 46053
rect 28634 46001 28686 46053
rect 28686 46001 28688 46053
rect 28632 45999 28688 46001
rect 28843 46053 28899 46055
rect 28843 46001 28845 46053
rect 28845 46001 28897 46053
rect 28897 46001 28899 46053
rect 28843 45999 28899 46001
rect 29054 46053 29110 46055
rect 29054 46001 29056 46053
rect 29056 46001 29108 46053
rect 29108 46001 29110 46053
rect 29054 45999 29110 46001
rect 56013 46053 56069 46055
rect 56013 46001 56015 46053
rect 56015 46001 56067 46053
rect 56067 46001 56069 46053
rect 56013 45999 56069 46001
rect 56224 46053 56280 46055
rect 56224 46001 56226 46053
rect 56226 46001 56278 46053
rect 56278 46001 56280 46053
rect 56224 45999 56280 46001
rect 56435 46053 56491 46055
rect 56435 46001 56437 46053
rect 56437 46001 56489 46053
rect 56489 46001 56491 46053
rect 56435 45999 56491 46001
rect 56646 46053 56702 46055
rect 56646 46001 56648 46053
rect 56648 46001 56700 46053
rect 56700 46001 56702 46053
rect 56646 45999 56702 46001
rect 56857 46053 56913 46055
rect 56857 46001 56859 46053
rect 56859 46001 56911 46053
rect 56911 46001 56913 46053
rect 56857 45999 56913 46001
rect 57068 46053 57124 46055
rect 57068 46001 57070 46053
rect 57070 46001 57122 46053
rect 57122 46001 57124 46053
rect 57068 45999 57124 46001
rect 57279 46053 57335 46055
rect 57279 46001 57281 46053
rect 57281 46001 57333 46053
rect 57333 46001 57335 46053
rect 57279 45999 57335 46001
rect 27788 44253 27844 44255
rect 27788 44201 27790 44253
rect 27790 44201 27842 44253
rect 27842 44201 27844 44253
rect 27788 44199 27844 44201
rect 27999 44253 28055 44255
rect 27999 44201 28001 44253
rect 28001 44201 28053 44253
rect 28053 44201 28055 44253
rect 27999 44199 28055 44201
rect 28210 44253 28266 44255
rect 28210 44201 28212 44253
rect 28212 44201 28264 44253
rect 28264 44201 28266 44253
rect 28210 44199 28266 44201
rect 28421 44253 28477 44255
rect 28421 44201 28423 44253
rect 28423 44201 28475 44253
rect 28475 44201 28477 44253
rect 28421 44199 28477 44201
rect 28632 44253 28688 44255
rect 28632 44201 28634 44253
rect 28634 44201 28686 44253
rect 28686 44201 28688 44253
rect 28632 44199 28688 44201
rect 28843 44253 28899 44255
rect 28843 44201 28845 44253
rect 28845 44201 28897 44253
rect 28897 44201 28899 44253
rect 28843 44199 28899 44201
rect 29054 44253 29110 44255
rect 29054 44201 29056 44253
rect 29056 44201 29108 44253
rect 29108 44201 29110 44253
rect 29054 44199 29110 44201
rect 56013 44253 56069 44255
rect 56013 44201 56015 44253
rect 56015 44201 56067 44253
rect 56067 44201 56069 44253
rect 56013 44199 56069 44201
rect 56224 44253 56280 44255
rect 56224 44201 56226 44253
rect 56226 44201 56278 44253
rect 56278 44201 56280 44253
rect 56224 44199 56280 44201
rect 56435 44253 56491 44255
rect 56435 44201 56437 44253
rect 56437 44201 56489 44253
rect 56489 44201 56491 44253
rect 56435 44199 56491 44201
rect 56646 44253 56702 44255
rect 56646 44201 56648 44253
rect 56648 44201 56700 44253
rect 56700 44201 56702 44253
rect 56646 44199 56702 44201
rect 56857 44253 56913 44255
rect 56857 44201 56859 44253
rect 56859 44201 56911 44253
rect 56911 44201 56913 44253
rect 56857 44199 56913 44201
rect 57068 44253 57124 44255
rect 57068 44201 57070 44253
rect 57070 44201 57122 44253
rect 57122 44201 57124 44253
rect 57068 44199 57124 44201
rect 57279 44253 57335 44255
rect 57279 44201 57281 44253
rect 57281 44201 57333 44253
rect 57333 44201 57335 44253
rect 57279 44199 57335 44201
rect 27788 42453 27844 42455
rect 27788 42401 27790 42453
rect 27790 42401 27842 42453
rect 27842 42401 27844 42453
rect 27788 42399 27844 42401
rect 27999 42453 28055 42455
rect 27999 42401 28001 42453
rect 28001 42401 28053 42453
rect 28053 42401 28055 42453
rect 27999 42399 28055 42401
rect 28210 42453 28266 42455
rect 28210 42401 28212 42453
rect 28212 42401 28264 42453
rect 28264 42401 28266 42453
rect 28210 42399 28266 42401
rect 28421 42453 28477 42455
rect 28421 42401 28423 42453
rect 28423 42401 28475 42453
rect 28475 42401 28477 42453
rect 28421 42399 28477 42401
rect 28632 42453 28688 42455
rect 28632 42401 28634 42453
rect 28634 42401 28686 42453
rect 28686 42401 28688 42453
rect 28632 42399 28688 42401
rect 28843 42453 28899 42455
rect 28843 42401 28845 42453
rect 28845 42401 28897 42453
rect 28897 42401 28899 42453
rect 28843 42399 28899 42401
rect 29054 42453 29110 42455
rect 29054 42401 29056 42453
rect 29056 42401 29108 42453
rect 29108 42401 29110 42453
rect 29054 42399 29110 42401
rect 56013 42453 56069 42455
rect 56013 42401 56015 42453
rect 56015 42401 56067 42453
rect 56067 42401 56069 42453
rect 56013 42399 56069 42401
rect 56224 42453 56280 42455
rect 56224 42401 56226 42453
rect 56226 42401 56278 42453
rect 56278 42401 56280 42453
rect 56224 42399 56280 42401
rect 56435 42453 56491 42455
rect 56435 42401 56437 42453
rect 56437 42401 56489 42453
rect 56489 42401 56491 42453
rect 56435 42399 56491 42401
rect 56646 42453 56702 42455
rect 56646 42401 56648 42453
rect 56648 42401 56700 42453
rect 56700 42401 56702 42453
rect 56646 42399 56702 42401
rect 56857 42453 56913 42455
rect 56857 42401 56859 42453
rect 56859 42401 56911 42453
rect 56911 42401 56913 42453
rect 56857 42399 56913 42401
rect 57068 42453 57124 42455
rect 57068 42401 57070 42453
rect 57070 42401 57122 42453
rect 57122 42401 57124 42453
rect 57068 42399 57124 42401
rect 57279 42453 57335 42455
rect 57279 42401 57281 42453
rect 57281 42401 57333 42453
rect 57333 42401 57335 42453
rect 57279 42399 57335 42401
rect 27788 40653 27844 40655
rect 27788 40601 27790 40653
rect 27790 40601 27842 40653
rect 27842 40601 27844 40653
rect 27788 40599 27844 40601
rect 27999 40653 28055 40655
rect 27999 40601 28001 40653
rect 28001 40601 28053 40653
rect 28053 40601 28055 40653
rect 27999 40599 28055 40601
rect 28210 40653 28266 40655
rect 28210 40601 28212 40653
rect 28212 40601 28264 40653
rect 28264 40601 28266 40653
rect 28210 40599 28266 40601
rect 28421 40653 28477 40655
rect 28421 40601 28423 40653
rect 28423 40601 28475 40653
rect 28475 40601 28477 40653
rect 28421 40599 28477 40601
rect 28632 40653 28688 40655
rect 28632 40601 28634 40653
rect 28634 40601 28686 40653
rect 28686 40601 28688 40653
rect 28632 40599 28688 40601
rect 28843 40653 28899 40655
rect 28843 40601 28845 40653
rect 28845 40601 28897 40653
rect 28897 40601 28899 40653
rect 28843 40599 28899 40601
rect 29054 40653 29110 40655
rect 29054 40601 29056 40653
rect 29056 40601 29108 40653
rect 29108 40601 29110 40653
rect 29054 40599 29110 40601
rect 56013 40653 56069 40655
rect 56013 40601 56015 40653
rect 56015 40601 56067 40653
rect 56067 40601 56069 40653
rect 56013 40599 56069 40601
rect 56224 40653 56280 40655
rect 56224 40601 56226 40653
rect 56226 40601 56278 40653
rect 56278 40601 56280 40653
rect 56224 40599 56280 40601
rect 56435 40653 56491 40655
rect 56435 40601 56437 40653
rect 56437 40601 56489 40653
rect 56489 40601 56491 40653
rect 56435 40599 56491 40601
rect 56646 40653 56702 40655
rect 56646 40601 56648 40653
rect 56648 40601 56700 40653
rect 56700 40601 56702 40653
rect 56646 40599 56702 40601
rect 56857 40653 56913 40655
rect 56857 40601 56859 40653
rect 56859 40601 56911 40653
rect 56911 40601 56913 40653
rect 56857 40599 56913 40601
rect 57068 40653 57124 40655
rect 57068 40601 57070 40653
rect 57070 40601 57122 40653
rect 57122 40601 57124 40653
rect 57068 40599 57124 40601
rect 57279 40653 57335 40655
rect 57279 40601 57281 40653
rect 57281 40601 57333 40653
rect 57333 40601 57335 40653
rect 57279 40599 57335 40601
rect 27788 38853 27844 38855
rect 27788 38801 27790 38853
rect 27790 38801 27842 38853
rect 27842 38801 27844 38853
rect 27788 38799 27844 38801
rect 27999 38853 28055 38855
rect 27999 38801 28001 38853
rect 28001 38801 28053 38853
rect 28053 38801 28055 38853
rect 27999 38799 28055 38801
rect 28210 38853 28266 38855
rect 28210 38801 28212 38853
rect 28212 38801 28264 38853
rect 28264 38801 28266 38853
rect 28210 38799 28266 38801
rect 28421 38853 28477 38855
rect 28421 38801 28423 38853
rect 28423 38801 28475 38853
rect 28475 38801 28477 38853
rect 28421 38799 28477 38801
rect 28632 38853 28688 38855
rect 28632 38801 28634 38853
rect 28634 38801 28686 38853
rect 28686 38801 28688 38853
rect 28632 38799 28688 38801
rect 28843 38853 28899 38855
rect 28843 38801 28845 38853
rect 28845 38801 28897 38853
rect 28897 38801 28899 38853
rect 28843 38799 28899 38801
rect 29054 38853 29110 38855
rect 29054 38801 29056 38853
rect 29056 38801 29108 38853
rect 29108 38801 29110 38853
rect 29054 38799 29110 38801
rect 56013 38853 56069 38855
rect 56013 38801 56015 38853
rect 56015 38801 56067 38853
rect 56067 38801 56069 38853
rect 56013 38799 56069 38801
rect 56224 38853 56280 38855
rect 56224 38801 56226 38853
rect 56226 38801 56278 38853
rect 56278 38801 56280 38853
rect 56224 38799 56280 38801
rect 56435 38853 56491 38855
rect 56435 38801 56437 38853
rect 56437 38801 56489 38853
rect 56489 38801 56491 38853
rect 56435 38799 56491 38801
rect 56646 38853 56702 38855
rect 56646 38801 56648 38853
rect 56648 38801 56700 38853
rect 56700 38801 56702 38853
rect 56646 38799 56702 38801
rect 56857 38853 56913 38855
rect 56857 38801 56859 38853
rect 56859 38801 56911 38853
rect 56911 38801 56913 38853
rect 56857 38799 56913 38801
rect 57068 38853 57124 38855
rect 57068 38801 57070 38853
rect 57070 38801 57122 38853
rect 57122 38801 57124 38853
rect 57068 38799 57124 38801
rect 57279 38853 57335 38855
rect 57279 38801 57281 38853
rect 57281 38801 57333 38853
rect 57333 38801 57335 38853
rect 57279 38799 57335 38801
rect 27788 37053 27844 37055
rect 27788 37001 27790 37053
rect 27790 37001 27842 37053
rect 27842 37001 27844 37053
rect 27788 36999 27844 37001
rect 27999 37053 28055 37055
rect 27999 37001 28001 37053
rect 28001 37001 28053 37053
rect 28053 37001 28055 37053
rect 27999 36999 28055 37001
rect 28210 37053 28266 37055
rect 28210 37001 28212 37053
rect 28212 37001 28264 37053
rect 28264 37001 28266 37053
rect 28210 36999 28266 37001
rect 28421 37053 28477 37055
rect 28421 37001 28423 37053
rect 28423 37001 28475 37053
rect 28475 37001 28477 37053
rect 28421 36999 28477 37001
rect 28632 37053 28688 37055
rect 28632 37001 28634 37053
rect 28634 37001 28686 37053
rect 28686 37001 28688 37053
rect 28632 36999 28688 37001
rect 28843 37053 28899 37055
rect 28843 37001 28845 37053
rect 28845 37001 28897 37053
rect 28897 37001 28899 37053
rect 28843 36999 28899 37001
rect 29054 37053 29110 37055
rect 29054 37001 29056 37053
rect 29056 37001 29108 37053
rect 29108 37001 29110 37053
rect 29054 36999 29110 37001
rect 56013 37053 56069 37055
rect 56013 37001 56015 37053
rect 56015 37001 56067 37053
rect 56067 37001 56069 37053
rect 56013 36999 56069 37001
rect 56224 37053 56280 37055
rect 56224 37001 56226 37053
rect 56226 37001 56278 37053
rect 56278 37001 56280 37053
rect 56224 36999 56280 37001
rect 56435 37053 56491 37055
rect 56435 37001 56437 37053
rect 56437 37001 56489 37053
rect 56489 37001 56491 37053
rect 56435 36999 56491 37001
rect 56646 37053 56702 37055
rect 56646 37001 56648 37053
rect 56648 37001 56700 37053
rect 56700 37001 56702 37053
rect 56646 36999 56702 37001
rect 56857 37053 56913 37055
rect 56857 37001 56859 37053
rect 56859 37001 56911 37053
rect 56911 37001 56913 37053
rect 56857 36999 56913 37001
rect 57068 37053 57124 37055
rect 57068 37001 57070 37053
rect 57070 37001 57122 37053
rect 57122 37001 57124 37053
rect 57068 36999 57124 37001
rect 57279 37053 57335 37055
rect 57279 37001 57281 37053
rect 57281 37001 57333 37053
rect 57333 37001 57335 37053
rect 57279 36999 57335 37001
rect 36958 35825 37014 35881
rect 37169 35825 37225 35881
rect 37381 35825 37437 35881
rect 37592 35825 37648 35881
rect 27474 26743 27530 26799
rect 27686 26743 27742 26799
rect 27474 26525 27530 26581
rect 27686 26525 27742 26581
rect 26450 26126 26610 26286
rect 26092 25807 26252 25967
rect 25756 25487 25916 25647
rect 25421 25168 25581 25328
rect 25081 24477 25241 24637
rect 24744 24156 24904 24316
rect 24416 23835 24576 23995
rect 24057 23513 24217 23673
rect 27474 24972 27530 25028
rect 27686 24972 27742 25028
rect 27474 24754 27530 24810
rect 27686 24754 27742 24810
rect 26924 20410 27084 20570
rect 26924 20066 27084 20226
rect 26465 19532 26625 19692
rect 26107 19187 26267 19347
rect 25771 18867 25931 19027
rect 25434 18524 25594 18684
rect 25094 18190 25254 18350
rect 24757 17817 24917 17977
rect 24429 17496 24589 17656
rect 24069 17157 24229 17317
rect 57381 26743 57437 26799
rect 57593 26743 57649 26799
rect 57381 26525 57437 26581
rect 57593 26525 57649 26581
rect 51766 9811 51822 9971
rect 49906 8900 50066 8956
rect 27474 7479 27530 7535
rect 27686 7479 27742 7535
rect 27474 7261 27530 7317
rect 27686 7261 27742 7317
rect 27474 7043 27530 7099
rect 27686 7043 27742 7099
rect 27474 6064 27530 6120
rect 27686 6064 27742 6120
rect 27474 5846 27530 5902
rect 27686 5846 27742 5902
rect 26859 5483 26915 5539
rect 27071 5483 27127 5539
rect 26859 5265 26915 5321
rect 27071 5265 27127 5321
rect 26859 4472 26915 4528
rect 27071 4472 27127 4528
rect 26859 4254 26915 4310
rect 27071 4254 27127 4310
rect 57381 6064 57437 6120
rect 57593 6064 57649 6120
rect 57381 5846 57437 5902
rect 57593 5846 57649 5902
rect 27474 3781 27530 3837
rect 27686 3781 27742 3837
rect 27474 3563 27530 3619
rect 27686 3563 27742 3619
rect 28801 3781 28857 3837
rect 28801 3563 28857 3619
rect 43800 2988 43960 3044
rect 57381 3781 57437 3837
rect 57593 3781 57649 3837
rect 57381 3563 57437 3619
rect 57593 3563 57649 3619
rect 57996 32032 58052 32088
rect 58208 32032 58264 32088
rect 57996 31814 58052 31870
rect 58208 31814 58264 31870
rect 57996 31596 58052 31652
rect 58208 31596 58264 31652
rect 58048 20410 58208 20570
rect 58048 20066 58208 20226
rect 57996 5483 58052 5539
rect 58208 5483 58264 5539
rect 57996 5265 58052 5321
rect 58208 5265 58264 5321
rect 57996 4472 58052 4528
rect 58208 4472 58264 4528
rect 57996 4254 58052 4310
rect 58208 4254 58264 4310
<< metal3 >>
rect 1401 52976 2401 53776
rect 2626 53168 3626 53776
rect 4137 52976 5137 53776
rect 5362 53168 6362 53776
rect 6801 52976 7801 53776
rect 8026 53168 9026 53776
rect 9537 52976 10537 53776
rect 10762 53168 11762 53776
rect 12201 52976 13201 53776
rect 13426 53168 14426 53776
rect 14937 52976 15937 53776
rect 16162 53168 17162 53776
rect 17601 52976 18601 53776
rect 18826 53168 19826 53776
rect 20653 52976 21653 53776
rect 22258 53168 23258 53776
rect 23483 52976 24483 53776
rect 25158 53168 26158 53776
rect 26572 52976 27572 53776
rect 27877 53168 28877 53776
rect 29273 53168 30273 53776
rect 30710 52976 31710 53776
rect 32381 53168 33381 53776
rect 34024 53168 35024 53776
rect 35415 52976 36415 53776
rect 36948 53168 37948 53776
rect 38585 52976 39585 53776
rect 39882 53168 40882 53776
rect 41230 52976 42230 53776
rect 42430 53168 43430 53776
rect 43713 53168 44713 53776
rect 45069 52976 46069 53776
rect 46313 52976 47313 53776
rect 47538 53168 48538 53776
rect 48901 52976 49901 53776
rect 50465 53168 51465 53776
rect 52569 52976 53569 53776
rect 54262 52976 55262 53776
rect 55990 53168 56990 53776
rect 57547 52976 58547 53776
rect 58791 53168 59791 53776
rect 60977 52976 61977 53776
rect 62202 53168 63202 53776
rect 63713 52976 64713 53776
rect 64938 53168 65938 53776
rect 66377 52976 67377 53776
rect 67602 53168 68602 53776
rect 69113 52976 70113 53776
rect 70338 53168 71338 53776
rect 71777 52976 72777 53776
rect 73002 53168 74002 53776
rect 74513 52976 75513 53776
rect 75738 53168 76738 53776
rect 77177 52976 78177 53776
rect 78402 53168 79402 53776
rect 80229 52976 81229 53776
rect 81834 53168 82834 53776
rect 83059 52976 84059 53776
rect 84666 52976 85666 53776
rect 0 51976 86372 52976
rect 0 51626 1014 51776
rect 0 51528 27779 51626
rect 58791 51576 59517 51591
rect 85358 51576 86372 51776
rect 58791 51528 86372 51576
rect 0 51455 86372 51528
rect 0 51399 27788 51455
rect 27844 51399 27999 51455
rect 28055 51399 28210 51455
rect 28266 51399 28421 51455
rect 28477 51399 28632 51455
rect 28688 51399 28843 51455
rect 28899 51399 29054 51455
rect 29110 51399 56013 51455
rect 56069 51399 56224 51455
rect 56280 51399 56435 51455
rect 56491 51399 56646 51455
rect 56702 51399 56857 51455
rect 56913 51399 57068 51455
rect 57124 51399 57279 51455
rect 57335 51399 86372 51455
rect 0 51327 86372 51399
rect 0 51226 27779 51327
rect 30402 51326 54622 51327
rect 58791 51276 86372 51327
rect 58791 51258 59517 51276
rect 0 51076 1014 51226
rect 85358 51076 86372 51276
rect 0 50176 1706 50876
rect 56271 50866 61644 51068
rect 41865 50613 42045 50623
rect 41865 50453 41875 50613
rect 42035 50453 42045 50613
rect 41865 50443 42045 50453
rect 84666 50176 86372 50876
rect 0 49776 1014 49976
rect 85358 49776 86372 49976
rect 0 49726 27272 49776
rect 30403 49726 54622 49728
rect 59421 49726 86372 49776
rect 0 49655 86372 49726
rect 0 49599 27788 49655
rect 27844 49599 27999 49655
rect 28055 49599 28210 49655
rect 28266 49599 28421 49655
rect 28477 49599 28632 49655
rect 28688 49599 28843 49655
rect 28899 49599 29054 49655
rect 29110 49599 56013 49655
rect 56069 49599 56224 49655
rect 56280 49599 56435 49655
rect 56491 49599 56646 49655
rect 56702 49599 56857 49655
rect 56913 49599 57068 49655
rect 57124 49599 57279 49655
rect 57335 49599 86372 49655
rect 0 49526 86372 49599
rect 0 49476 27272 49526
rect 59421 49476 86372 49526
rect 0 49276 1014 49476
rect 85358 49276 86372 49476
rect 0 48376 1706 49076
rect 84666 48376 86372 49076
rect 0 47976 1014 48176
rect 85358 47976 86372 48176
rect 0 47926 27272 47976
rect 30403 47926 54622 47928
rect 59421 47926 86372 47976
rect 0 47855 86372 47926
rect 0 47799 27788 47855
rect 27844 47799 27999 47855
rect 28055 47799 28210 47855
rect 28266 47799 28421 47855
rect 28477 47799 28632 47855
rect 28688 47799 28843 47855
rect 28899 47799 29054 47855
rect 29110 47799 56013 47855
rect 56069 47799 56224 47855
rect 56280 47799 56435 47855
rect 56491 47799 56646 47855
rect 56702 47799 56857 47855
rect 56913 47799 57068 47855
rect 57124 47799 57279 47855
rect 57335 47799 86372 47855
rect 0 47726 86372 47799
rect 0 47676 27272 47726
rect 59421 47676 86372 47726
rect 0 47476 1014 47676
rect 85358 47476 86372 47676
rect 0 46576 1706 47276
rect 84666 46576 86372 47276
rect 0 46176 1014 46376
rect 85358 46176 86372 46376
rect 0 46126 27272 46176
rect 30403 46126 54622 46128
rect 59421 46126 86372 46176
rect 0 46055 86372 46126
rect 0 45999 27788 46055
rect 27844 45999 27999 46055
rect 28055 45999 28210 46055
rect 28266 45999 28421 46055
rect 28477 45999 28632 46055
rect 28688 45999 28843 46055
rect 28899 45999 29054 46055
rect 29110 45999 56013 46055
rect 56069 45999 56224 46055
rect 56280 45999 56435 46055
rect 56491 45999 56646 46055
rect 56702 45999 56857 46055
rect 56913 45999 57068 46055
rect 57124 45999 57279 46055
rect 57335 45999 86372 46055
rect 0 45926 86372 45999
rect 0 45876 27272 45926
rect 59421 45876 86372 45926
rect 0 45676 1014 45876
rect 85358 45676 86372 45876
rect 0 44776 1706 45476
rect 84666 44776 86372 45476
rect 0 44376 1014 44576
rect 85358 44376 86372 44576
rect 0 44326 27272 44376
rect 30403 44326 54622 44328
rect 59421 44326 86372 44376
rect 0 44255 86372 44326
rect 0 44199 27788 44255
rect 27844 44199 27999 44255
rect 28055 44199 28210 44255
rect 28266 44199 28421 44255
rect 28477 44199 28632 44255
rect 28688 44199 28843 44255
rect 28899 44199 29054 44255
rect 29110 44199 56013 44255
rect 56069 44199 56224 44255
rect 56280 44199 56435 44255
rect 56491 44199 56646 44255
rect 56702 44199 56857 44255
rect 56913 44199 57068 44255
rect 57124 44199 57279 44255
rect 57335 44199 86372 44255
rect 0 44126 86372 44199
rect 0 44076 27272 44126
rect 59421 44076 86372 44126
rect 0 43876 1014 44076
rect 85358 43876 86372 44076
rect 0 42976 1706 43676
rect 84666 42976 86372 43676
rect 0 42576 1014 42776
rect 85358 42576 86372 42776
rect 0 42526 27272 42576
rect 30403 42526 54622 42528
rect 59421 42526 86372 42576
rect 0 42455 86372 42526
rect 0 42399 27788 42455
rect 27844 42399 27999 42455
rect 28055 42399 28210 42455
rect 28266 42399 28421 42455
rect 28477 42399 28632 42455
rect 28688 42399 28843 42455
rect 28899 42399 29054 42455
rect 29110 42399 56013 42455
rect 56069 42399 56224 42455
rect 56280 42399 56435 42455
rect 56491 42399 56646 42455
rect 56702 42399 56857 42455
rect 56913 42399 57068 42455
rect 57124 42399 57279 42455
rect 57335 42399 86372 42455
rect 0 42326 86372 42399
rect 0 42276 27272 42326
rect 59421 42276 86372 42326
rect 0 42076 1014 42276
rect 85358 42076 86372 42276
rect 0 41176 1706 41876
rect 84666 41176 86372 41876
rect 0 40776 1014 40976
rect 85358 40776 86372 40976
rect 0 40726 27272 40776
rect 30403 40726 54622 40728
rect 59421 40726 86372 40776
rect 0 40655 86372 40726
rect 0 40599 27788 40655
rect 27844 40599 27999 40655
rect 28055 40599 28210 40655
rect 28266 40599 28421 40655
rect 28477 40599 28632 40655
rect 28688 40599 28843 40655
rect 28899 40599 29054 40655
rect 29110 40599 56013 40655
rect 56069 40599 56224 40655
rect 56280 40599 56435 40655
rect 56491 40599 56646 40655
rect 56702 40599 56857 40655
rect 56913 40599 57068 40655
rect 57124 40599 57279 40655
rect 57335 40599 86372 40655
rect 0 40526 86372 40599
rect 0 40476 27272 40526
rect 59421 40476 86372 40526
rect 0 40276 1014 40476
rect 85358 40276 86372 40476
rect 0 39376 1706 40076
rect 84666 39376 86372 40076
rect 0 38976 1014 39176
rect 85358 38976 86372 39176
rect 0 38926 27272 38976
rect 30403 38926 54622 38928
rect 59421 38926 86372 38976
rect 0 38855 86372 38926
rect 0 38799 27788 38855
rect 27844 38799 27999 38855
rect 28055 38799 28210 38855
rect 28266 38799 28421 38855
rect 28477 38799 28632 38855
rect 28688 38799 28843 38855
rect 28899 38799 29054 38855
rect 29110 38799 56013 38855
rect 56069 38799 56224 38855
rect 56280 38799 56435 38855
rect 56491 38799 56646 38855
rect 56702 38799 56857 38855
rect 56913 38799 57068 38855
rect 57124 38799 57279 38855
rect 57335 38799 86372 38855
rect 0 38726 86372 38799
rect 0 38676 27272 38726
rect 59421 38676 86372 38726
rect 0 38476 1014 38676
rect 85358 38476 86372 38676
rect 0 37576 1706 38276
rect 84666 37576 86372 38276
rect 0 37176 1014 37376
rect 85358 37176 86372 37376
rect 0 37126 27272 37176
rect 30403 37126 54622 37128
rect 59421 37126 86372 37176
rect 0 37055 86372 37126
rect 0 36999 27788 37055
rect 27844 36999 27999 37055
rect 28055 36999 28210 37055
rect 28266 36999 28421 37055
rect 28477 36999 28632 37055
rect 28688 36999 28843 37055
rect 28899 36999 29054 37055
rect 29110 36999 56013 37055
rect 56069 36999 56224 37055
rect 56280 36999 56435 37055
rect 56491 36999 56646 37055
rect 56702 36999 56857 37055
rect 56913 36999 57068 37055
rect 57124 36999 57279 37055
rect 57335 36999 86372 37055
rect 0 36926 86372 36999
rect 0 36876 27272 36926
rect 59421 36876 86372 36926
rect 0 36676 1014 36876
rect 85358 36676 86372 36876
rect 0 35776 1706 36476
rect 36863 35881 37743 35920
rect 36863 35825 36958 35881
rect 37014 35825 37169 35881
rect 37225 35825 37381 35881
rect 37437 35825 37592 35881
rect 37648 35825 37743 35881
rect 0 34536 27828 35326
rect 2095 34125 2188 34126
rect 0 34124 25085 34125
rect 0 32318 27214 34124
rect 36863 33927 37743 35825
rect 84666 35776 86372 36476
rect 57369 34536 86372 35326
rect 61853 34124 72383 34125
rect 72653 34124 86372 34125
rect 0 32316 25085 32318
rect 0 32315 3011 32316
rect 0 29714 1706 32315
rect 27387 32311 28929 33263
rect 56135 32311 57736 33263
rect 57908 32315 86372 34124
rect 57908 32199 58351 32315
rect 26772 32088 58351 32199
rect 26772 32032 26859 32088
rect 26915 32032 27071 32088
rect 27127 32032 57996 32088
rect 58052 32032 58208 32088
rect 58264 32032 58351 32088
rect 26772 31870 58351 32032
rect 26772 31814 26859 31870
rect 26915 31814 27071 31870
rect 27127 31814 57996 31870
rect 58052 31814 58208 31870
rect 58264 31814 58351 31870
rect 26772 31652 58351 31814
rect 26772 31596 26859 31652
rect 26915 31596 27071 31652
rect 27127 31596 57996 31652
rect 58052 31596 58208 31652
rect 58264 31596 58351 31652
rect 26772 31486 58351 31596
rect 25293 30443 28929 31352
rect 56186 30443 59524 31352
rect 26772 29714 58351 30105
rect 84666 29714 86372 32315
rect 0 29430 86372 29714
rect 0 26890 26070 28416
rect 26772 27382 58351 29430
rect 58785 26890 86372 28416
rect 0 26799 27828 26890
rect 0 26743 27474 26799
rect 27530 26743 27686 26799
rect 27742 26743 27828 26799
rect 0 26581 27828 26743
rect 0 26525 27474 26581
rect 27530 26525 27686 26581
rect 27742 26525 27828 26581
rect 0 26435 27828 26525
rect 57295 26799 86372 26890
rect 57295 26743 57381 26799
rect 57437 26743 57593 26799
rect 57649 26743 86372 26799
rect 57295 26581 86372 26743
rect 57295 26525 57381 26581
rect 57437 26525 57593 26581
rect 57649 26525 86372 26581
rect 57295 26435 86372 26525
rect 6921 26434 8163 26435
rect 17721 26434 18963 26435
rect 66497 26434 67739 26435
rect 77297 26434 78539 26435
rect 23828 26286 26642 26324
rect 23828 26126 26450 26286
rect 26610 26126 26642 26286
rect 23828 26109 26642 26126
rect 23828 25967 26285 26002
rect 23828 25807 26092 25967
rect 26252 25807 26285 25967
rect 23828 25787 26285 25807
rect 23828 25647 25949 25681
rect 23828 25487 25756 25647
rect 25916 25487 25949 25647
rect 23828 25466 25949 25487
rect 23828 25328 25614 25359
rect 23828 25168 25421 25328
rect 25581 25168 25614 25328
rect 23828 25144 25614 25168
rect 27382 25028 29699 25208
rect 27382 24972 27474 25028
rect 27530 24972 27686 25028
rect 27742 24972 29699 25028
rect 27382 24810 29699 24972
rect 27382 24754 27474 24810
rect 27530 24754 27686 24810
rect 27742 24754 29699 24810
rect 23828 24637 25274 24667
rect 23828 24477 25081 24637
rect 25241 24477 25274 24637
rect 27382 24526 29699 24754
rect 23828 24452 25274 24477
rect 23828 24316 24935 24345
rect 23828 24156 24744 24316
rect 24904 24156 24935 24316
rect 23828 24130 24935 24156
rect 23828 23995 24607 24024
rect 0 23380 1706 23938
rect 23828 23835 24416 23995
rect 24576 23835 24607 23995
rect 23828 23809 24607 23835
rect 24047 23673 24227 23683
rect 24047 23513 24057 23673
rect 24217 23513 24227 23673
rect 24047 23503 24227 23513
rect 26770 23380 58348 24278
rect 84666 23380 86372 23938
rect 0 23370 86372 23380
rect 0 22938 27214 23370
rect 27387 22291 57677 23199
rect 57908 22938 86372 23370
rect 57908 22937 83763 22938
rect 27387 22282 27826 22291
rect 0 21827 27826 22282
rect 0 21282 1014 21827
rect 24036 21826 27826 21827
rect 56078 22282 57677 22291
rect 56078 21827 86372 22282
rect 56078 21826 83763 21827
rect 44432 21707 55645 21708
rect 29521 21625 55645 21707
rect 29513 20739 55645 21625
rect 85358 21282 86372 21827
rect 0 20570 86372 20739
rect 0 20410 26924 20570
rect 27084 20410 58048 20570
rect 58208 20410 86372 20570
rect 0 20226 86372 20410
rect 0 20066 26924 20226
rect 27084 20066 58048 20226
rect 58208 20066 86372 20226
rect 0 19969 86372 20066
rect 0 18016 24250 19969
rect 26435 19692 29403 19731
rect 26435 19532 26465 19692
rect 26625 19532 29403 19692
rect 26435 19502 29403 19532
rect 55720 19502 58817 19731
rect 26077 19347 29403 19391
rect 26077 19187 26107 19347
rect 26267 19187 29403 19347
rect 26077 19162 29403 19187
rect 55720 19162 59177 19391
rect 25742 19027 29403 19051
rect 25742 18867 25771 19027
rect 25931 18867 29403 19027
rect 25742 18822 29403 18867
rect 55720 18822 59515 19051
rect 25406 18684 29403 18711
rect 25406 18524 25434 18684
rect 25594 18524 29403 18684
rect 25406 18482 29403 18524
rect 55720 18482 59846 18711
rect 25066 18350 29403 18371
rect 25066 18190 25094 18350
rect 25254 18190 29403 18350
rect 25066 18142 29403 18190
rect 55720 18142 60184 18371
rect 24730 17977 29403 18031
rect 24730 17817 24757 17977
rect 24917 17817 29403 17977
rect 24730 17802 29403 17817
rect 55720 17802 60525 18031
rect 61807 18016 86372 19969
rect 61825 18015 83763 18016
rect 0 16597 23678 17730
rect 24401 17656 29403 17691
rect 24401 17496 24429 17656
rect 24589 17496 29403 17656
rect 24401 17462 29403 17496
rect 55720 17462 60855 17691
rect 24042 17317 29403 17351
rect 24042 17157 24069 17317
rect 24229 17157 29403 17317
rect 24042 17122 29403 17157
rect 55720 17122 61205 17351
rect 61807 16784 86372 17730
rect 24111 16597 27828 16598
rect 0 15015 27828 16597
rect 46982 15015 86372 16784
rect 0 14968 86372 15015
rect 0 14966 55645 14968
rect 0 14936 51760 14966
rect 0 14491 47683 14936
rect 0 14329 45977 14491
rect 0 14328 24250 14329
rect 24047 14178 27214 14179
rect 0 13461 27214 14178
rect 0 12846 1706 13461
rect 24047 12934 27214 13461
rect 27387 13760 45977 14329
rect 57295 14328 86372 14968
rect 57295 14327 83763 14328
rect 83169 14178 84221 14179
rect 61807 14177 72429 14178
rect 72607 14177 86372 14178
rect 59826 13866 60026 14017
rect 61773 13866 86372 14177
rect 27387 13245 49775 13760
rect 29478 13243 49775 13245
rect 41493 13078 49775 13243
rect 50228 13461 86372 13866
rect 24047 12847 34761 12934
rect 23821 12846 34761 12847
rect 0 12574 34761 12846
rect 50228 12846 58421 13461
rect 59826 12846 60026 13461
rect 83169 12846 84221 12847
rect 84666 12846 86372 13461
rect 50228 12574 86372 12846
rect 0 12046 86372 12574
rect 0 12036 24250 12046
rect 26772 12036 86372 12046
rect 26772 12035 84999 12036
rect 26772 11844 58351 12035
rect 29478 11697 58351 11844
rect 0 11491 3011 11493
rect 24047 11491 27828 11493
rect 0 10176 27828 11491
rect 29478 10756 41516 11697
rect 2229 10175 24250 10176
rect 2249 10174 24250 10175
rect 23612 9942 29221 10030
rect 34741 9972 41516 10756
rect 42261 11491 57736 11527
rect 61825 11491 86372 11493
rect 42261 10740 86372 11491
rect 24047 9515 28729 9516
rect 0 8154 28729 9515
rect 29133 9302 29221 9942
rect 41857 9502 51430 10420
rect 51750 10097 54952 10185
rect 57295 10176 86372 10740
rect 61805 10175 84482 10176
rect 61825 10173 84482 10175
rect 51750 9971 51838 10097
rect 51750 9811 51766 9971
rect 51822 9811 51838 9971
rect 54864 10028 54952 10097
rect 54864 9940 62145 10028
rect 51750 9801 51838 9811
rect 58688 9681 61743 9777
rect 57909 9514 62278 9516
rect 83361 9514 86372 9515
rect 29133 9214 41656 9302
rect 41568 8972 41656 9214
rect 41857 9165 55482 9502
rect 41568 8956 50076 8972
rect 41568 8900 49906 8956
rect 50066 8900 50076 8956
rect 41568 8884 50076 8900
rect 50922 8888 55482 9165
rect 0 8153 24250 8154
rect 0 8152 3011 8153
rect 28178 7652 28729 8154
rect 29513 7900 41397 8582
rect 0 7595 3011 7596
rect 23625 7595 27828 7596
rect 0 7535 27828 7595
rect 0 7479 27474 7535
rect 27530 7479 27686 7535
rect 27742 7479 27828 7535
rect 0 7317 27828 7479
rect 0 7261 27474 7317
rect 27530 7261 27686 7317
rect 27742 7261 27828 7317
rect 0 7099 27828 7261
rect 0 7043 27474 7099
rect 27530 7043 27686 7099
rect 27742 7043 27828 7099
rect 28178 7084 34622 7652
rect 0 6982 27828 7043
rect 0 6199 1014 6982
rect 2226 6981 24250 6982
rect 2249 6980 24250 6981
rect 23625 6306 29058 6875
rect 29537 6744 34622 7084
rect 34860 7392 41397 7900
rect 50922 7596 57736 8888
rect 57909 8154 86372 9514
rect 61802 8153 86372 8154
rect 61825 8152 86372 8153
rect 50922 7595 62747 7596
rect 83361 7595 86372 7596
rect 50922 7392 86372 7595
rect 34860 6984 86372 7392
rect 34860 6592 55482 6984
rect 57295 6982 86372 6984
rect 61802 6981 84787 6982
rect 61825 6980 84787 6981
rect 34860 6573 41397 6592
rect 29458 6199 41397 6573
rect 0 6198 3011 6199
rect 23687 6198 41397 6199
rect 0 6177 41397 6198
rect 50922 6199 55482 6592
rect 56065 6306 62747 6875
rect 85358 6199 86372 6982
rect 50922 6198 62429 6199
rect 83361 6198 86372 6199
rect 0 6120 34622 6177
rect 0 6064 27474 6120
rect 27530 6064 27686 6120
rect 27742 6064 34622 6120
rect 0 5902 34622 6064
rect 0 5846 27474 5902
rect 27530 5846 27686 5902
rect 27742 5846 34622 5902
rect 0 5766 34622 5846
rect 29458 5665 34622 5766
rect 50922 6120 86372 6198
rect 50922 6064 57381 6120
rect 57437 6064 57593 6120
rect 57649 6064 86372 6120
rect 50922 5902 86372 6064
rect 50922 5846 57381 5902
rect 57437 5846 57593 5902
rect 57649 5846 86372 5902
rect 50922 5766 86372 5846
rect 23687 5629 27214 5630
rect 0 5539 27214 5629
rect 50922 5605 55482 5766
rect 57909 5629 62429 5630
rect 0 5483 26859 5539
rect 26915 5483 27071 5539
rect 27127 5483 27214 5539
rect 0 5321 27214 5483
rect 0 5265 26859 5321
rect 26915 5265 27071 5321
rect 27127 5265 27214 5321
rect 0 5175 27214 5265
rect 57909 5539 86372 5629
rect 57909 5483 57996 5539
rect 58052 5483 58208 5539
rect 58264 5483 86372 5539
rect 57909 5321 86372 5483
rect 57909 5265 57996 5321
rect 58052 5265 58208 5321
rect 58264 5265 86372 5321
rect 57909 5175 86372 5265
rect 0 5174 24250 5175
rect 61802 5174 86372 5175
rect 0 5173 3011 5174
rect 83361 5173 86372 5174
rect 0 4515 1712 5173
rect 57909 4619 62429 4621
rect 23909 4528 62429 4619
rect 23909 4515 26859 4528
rect 0 4472 26859 4515
rect 26915 4472 27071 4528
rect 27127 4472 57996 4528
rect 58052 4472 58208 4528
rect 58264 4515 62429 4528
rect 84660 4515 86372 5173
rect 58264 4472 86372 4515
rect 0 4310 86372 4472
rect 0 4254 26859 4310
rect 26915 4254 27071 4310
rect 27127 4254 57996 4310
rect 58052 4254 58208 4310
rect 58264 4254 86372 4310
rect 0 4166 86372 4254
rect 0 4164 59323 4166
rect 0 4060 24341 4164
rect 61788 4060 86372 4166
rect 27438 3875 27778 3876
rect 28764 3875 28894 3876
rect 41774 3875 41904 3876
rect 42299 3875 42429 3876
rect 46873 3875 47003 3876
rect 47321 3875 47451 3876
rect 47769 3875 47899 3876
rect 48217 3875 48347 3876
rect 57345 3875 61215 3876
rect 23909 3837 61215 3875
rect 23909 3781 27474 3837
rect 27530 3781 27686 3837
rect 27742 3781 28801 3837
rect 28857 3781 57381 3837
rect 57437 3781 57593 3837
rect 57649 3781 61215 3837
rect 23909 3772 61215 3781
rect 0 3619 86372 3772
rect 0 3563 27474 3619
rect 27530 3563 27686 3619
rect 27742 3563 28801 3619
rect 28857 3563 57381 3619
rect 57437 3563 57593 3619
rect 57649 3563 86372 3619
rect 0 3524 86372 3563
rect 0 3421 24341 3524
rect 0 3420 3011 3421
rect 60886 3420 86372 3524
rect 0 2854 1000 3420
rect 24169 3044 62588 3066
rect 24169 2988 43800 3044
rect 43960 2988 62588 3044
rect 24169 2978 62588 2988
rect 85358 2854 86372 3420
rect 0 2502 86372 2854
rect 0 1232 86372 2232
rect 706 0 1706 1232
rect 2039 0 3039 1232
rect 3442 0 4442 1232
rect 4642 0 5642 932
rect 5842 0 6842 1232
rect 7042 0 8042 1232
rect 8242 0 9242 1232
rect 9442 0 10442 932
rect 10642 0 11642 1232
rect 12443 0 13443 1232
rect 14242 0 15242 1232
rect 15442 0 16442 932
rect 16642 0 17642 1232
rect 17842 0 18842 1232
rect 19042 0 20042 1232
rect 20242 0 21242 932
rect 21910 0 22910 1232
rect 23110 0 24110 1232
rect 24410 0 25410 1232
rect 25710 0 26710 1232
rect 27010 0 28010 1232
rect 28310 0 29310 1232
rect 29610 0 30610 1232
rect 31324 0 32324 932
rect 33022 0 34022 932
rect 34831 0 35831 932
rect 36031 0 37031 1232
rect 38028 0 39028 932
rect 39228 0 40228 1232
rect 41233 0 42233 932
rect 42433 0 43433 1232
rect 43633 0 44633 932
rect 44833 0 45833 1232
rect 46033 0 47033 932
rect 47233 0 48233 1232
rect 48566 0 49566 1232
rect 49876 0 50876 1232
rect 51233 0 52233 932
rect 52478 0 53478 932
rect 54458 0 55458 1232
rect 55758 0 56758 1232
rect 57058 0 58058 1232
rect 58358 0 59358 1232
rect 59658 0 60658 1232
rect 60958 0 61958 1232
rect 62295 0 63295 1232
rect 64218 0 65218 932
rect 65418 0 66418 1232
rect 66618 0 67618 1232
rect 67818 0 68818 1232
rect 69018 0 70018 932
rect 70218 0 71218 1232
rect 72017 0 73017 1232
rect 73818 0 74818 1232
rect 75018 0 76018 932
rect 76218 0 77218 1232
rect 77418 0 78418 1232
rect 78618 0 79618 1232
rect 79818 0 80818 932
rect 81018 0 82018 1232
rect 82419 0 83419 1232
rect 84666 0 85666 1232
use 128x8M8WM1_PWR_128x8m81  128x8M8WM1_PWR_128x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 1912 6592 83548 35222
use GF018_128x8M8WM1_lef_128x8m81  GF018_128x8M8WM1_lef_128x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 0
box 0 0 86372 53776
use G_ring_128x8m81  G_ring_128x8m81_0
timestamp 1666464484
transform 1 0 282 0 1 0
box 0 0 85816 53502
use M1_PSUB431059054877_128x8m81  M1_PSUB431059054877_128x8m81_0
timestamp 1666464484
transform 1 0 53710 0 1 2781
box -2884 -1144 2884 1144
use M1_PSUB4310590548712_128x8m81  M1_PSUB4310590548712_128x8m81_0
timestamp 1666464484
transform 1 0 34404 0 1 2781
box -5784 -1144 5784 1144
use M1_PSUB4310590548715_128x8m81  M1_PSUB4310590548715_128x8m81_0
timestamp 1666464484
transform 1 0 57403 0 1 1140
box -42 -42 242 51842
use M1_PSUB4310590548715_128x8m81  M1_PSUB4310590548715_128x8m81_1
timestamp 1666464484
transform 1 0 27521 0 1 1140
box -42 -42 242 51842
use M1_PSUB4310590548716_128x8m81  M1_PSUB4310590548716_128x8m81_0
timestamp 1666464484
transform 1 0 27869 0 1 34279
box -42 -42 29442 342
use M1_PSUB4310590548717_128x8m81  M1_PSUB4310590548717_128x8m81_0
timestamp 1666464484
transform 1 0 27869 0 1 36019
box -42 -42 642 16942
use M1_PSUB4310590548717_128x8m81  M1_PSUB4310590548717_128x8m81_1
timestamp 1666464484
transform 1 0 56655 0 1 36019
box -42 -42 642 16942
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_0
timestamp 1666464484
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_1
timestamp 1666464484
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_2
timestamp 1666464484
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_3
timestamp 1666464484
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_4
timestamp 1666464484
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_5
timestamp 1666464484
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_6
timestamp 1666464484
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_7
timestamp 1666464484
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_8
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_9
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_10
timestamp 1666464484
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_11
timestamp 1666464484
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_12
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_13
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_14
timestamp 1666464484
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_15
timestamp 1666464484
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_16
timestamp 1666464484
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_17
timestamp 1666464484
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_18
timestamp 1666464484
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M2_M1$$199747628_128x8m81  M2_M1$$199747628_128x8m81_19
timestamp 1666464484
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201260076_128x8m81  M2_M1$$201260076_128x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 19369
box -170 -14104 170 14104
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 4126
box -170 -502 170 502
use M2_M1$$201261100_128x8m81  M2_M1$$201261100_128x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 4126
box -170 -502 170 502
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_0
timestamp 1666464484
transform 1 0 82808 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_1
timestamp 1666464484
transform 1 0 51732 0 1 5173
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_2
timestamp 1666464484
transform 1 0 72743 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_3
timestamp 1666464484
transform 1 0 72293 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_4
timestamp 1666464484
transform 1 0 62228 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_5
timestamp 1666464484
transform 1 0 49986 0 1 6323
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_6
timestamp 1666464484
transform 1 0 40700 0 1 4878
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_7
timestamp 1666464484
transform 1 0 23517 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_8
timestamp 1666464484
transform 1 0 13167 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_9
timestamp 1666464484
transform 1 0 12717 0 1 1663
box 0 0 1 1
use M2_M1431059054870_128x8m81  M2_M1431059054870_128x8m81_10
timestamp 1666464484
transform 1 0 2652 0 1 1663
box 0 0 1 1
use M2_M1431059054873_128x8m81  M2_M1431059054873_128x8m81_0
timestamp 1666464484
transform 1 0 27590 0 1 34937
box -162 -348 162 348
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1666464484
transform 1 0 60601 0 1 35416
box 0 0 1 1
use M2_M14310590548711_128x8m81  M2_M14310590548711_128x8m81_0
timestamp 1666464484
transform 1 0 57507 0 1 34906
box -100 -348 100 348
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_0
timestamp 1666464484
transform 1 0 29818 0 1 785
box 0 0 1 1
use M2_M14310590548713_128x8m81  M2_M14310590548713_128x8m81_1
timestamp 1666464484
transform 1 0 29116 0 1 785
box 0 0 1 1
use M2_M14310590548719_128x8m81  M2_M14310590548719_128x8m81_0
timestamp 1666464484
transform 1 0 25674 0 1 51429
box -286 -162 286 162
use M2_M14310590548719_128x8m81  M2_M14310590548719_128x8m81_1
timestamp 1666464484
transform 1 0 59152 0 1 51429
box -286 -162 286 162
use M2_M14310590548721_128x8m81  M2_M14310590548721_128x8m81_0
timestamp 1666464484
transform 1 0 48818 0 1 764
box -162 -472 162 472
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 12783
box -170 -1046 170 1046
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 15671
box -170 -1046 170 1046
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 15463
box -170 -1046 170 1046
use M3_M2$$201248812_128x8m81  M3_M2$$201248812_128x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 13112
box -170 -1046 170 1046
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_0
timestamp 1666464484
transform -1 0 57515 0 1 10834
box -170 -611 170 611
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 8835
box -170 -611 170 611
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_2
timestamp 1666464484
transform 1 0 27608 0 1 10834
box -170 -611 170 611
use M3_M2$$201249836_128x8m81  M3_M2$$201249836_128x8m81_3
timestamp 1666464484
transform 1 0 26993 0 1 8835
box -170 -611 170 611
use M3_M2$$201250860_128x8m81  M3_M2$$201250860_128x8m81_0
timestamp 1666464484
transform -1 0 56505 0 1 6590
box -381 -284 381 284
use M3_M2$$201250860_128x8m81  M3_M2$$201250860_128x8m81_1
timestamp 1666464484
transform 1 0 28618 0 1 6590
box -381 -284 381 284
use M3_M2$$201251884_128x8m81  M3_M2$$201251884_128x8m81_0
timestamp 1666464484
transform 1 0 37303 0 1 35853
box 0 0 1 1
use M3_M2$$201252908_128x8m81  M3_M2$$201252908_128x8m81_0
timestamp 1666464484
transform 1 0 28829 0 1 3700
box 0 0 1 1
use M3_M2$$201253932_128x8m81  M3_M2$$201253932_128x8m81_0
timestamp 1666464484
transform 1 0 57515 0 1 8156
box -170 -1155 170 716
use M3_M2$$201254956_128x8m81  M3_M2$$201254956_128x8m81_0
timestamp 1666464484
transform 1 0 27608 0 1 13768
box -170 -502 170 502
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_0
timestamp 1666464484
transform 1 0 28449 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_1
timestamp 1666464484
transform 1 0 28449 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_2
timestamp 1666464484
transform 1 0 28449 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_3
timestamp 1666464484
transform 1 0 28449 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_4
timestamp 1666464484
transform 1 0 28449 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_5
timestamp 1666464484
transform 1 0 28449 0 1 37027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_6
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_7
timestamp 1666464484
transform 1 0 28449 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_8
timestamp 1666464484
transform 1 0 28449 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_9
timestamp 1666464484
transform 1 0 28449 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_10
timestamp 1666464484
transform 1 0 56674 0 1 38827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_11
timestamp 1666464484
transform 1 0 56674 0 1 40627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_12
timestamp 1666464484
transform 1 0 56674 0 1 42427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_13
timestamp 1666464484
transform 1 0 56674 0 1 44227
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_14
timestamp 1666464484
transform 1 0 56674 0 1 46027
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_15
timestamp 1666464484
transform 1 0 56674 0 1 47827
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_16
timestamp 1666464484
transform 1 0 56674 0 1 49627
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_17
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_18
timestamp 1666464484
transform 1 0 56674 0 1 51427
box 0 0 1 1
use M3_M2$$201258028_128x8m81  M3_M2$$201258028_128x8m81_19
timestamp 1666464484
transform 1 0 56674 0 1 37027
box 0 0 1 1
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_0
timestamp 1666464484
transform 1 0 27608 0 1 32786
box -170 -393 170 393
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_1
timestamp 1666464484
transform 1 0 27608 0 1 30897
box -170 -393 170 393
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_2
timestamp 1666464484
transform -1 0 57515 0 1 30897
box -170 -393 170 393
use M3_M2$$201412652_128x8m81  M3_M2$$201412652_128x8m81_3
timestamp 1666464484
transform -1 0 57515 0 1 32786
box -170 -393 170 393
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_0
timestamp 1666464484
transform 1 0 27608 0 1 7289
box 0 0 1 1
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_1
timestamp 1666464484
transform 1 0 26993 0 1 31842
box 0 0 1 1
use M3_M2$$201413676_128x8m81  M3_M2$$201413676_128x8m81_2
timestamp 1666464484
transform -1 0 58130 0 1 31842
box 0 0 1 1
use M3_M2$$201414700_128x8m81  M3_M2$$201414700_128x8m81_0
timestamp 1666464484
transform 1 0 26993 0 1 33221
box -170 -828 170 828
use M3_M2$$201414700_128x8m81  M3_M2$$201414700_128x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 33221
box -170 -828 170 828
use M3_M2$$201415724_128x8m81  M3_M2$$201415724_128x8m81_0
timestamp 1666464484
transform 1 0 26993 0 1 28743
box -170 -1264 170 1264
use M3_M2$$201415724_128x8m81  M3_M2$$201415724_128x8m81_1
timestamp 1666464484
transform -1 0 58130 0 1 28743
box -170 -1264 170 1264
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_0
timestamp 1666464484
transform -1 0 58130 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_1
timestamp 1666464484
transform -1 0 57515 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_2
timestamp 1666464484
transform -1 0 57515 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_3
timestamp 1666464484
transform -1 0 58130 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_4
timestamp 1666464484
transform -1 0 57515 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_5
timestamp 1666464484
transform 1 0 27608 0 1 3700
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_6
timestamp 1666464484
transform 1 0 26993 0 1 4391
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_7
timestamp 1666464484
transform 1 0 27608 0 1 5983
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_8
timestamp 1666464484
transform 1 0 26993 0 1 5402
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_9
timestamp 1666464484
transform 1 0 27608 0 1 26662
box 0 0 1 1
use M3_M2$$201416748_128x8m81  M3_M2$$201416748_128x8m81_10
timestamp 1666464484
transform 1 0 27608 0 1 24891
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1666464484
transform 0 -1 49986 1 0 8928
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_1
timestamp 1666464484
transform 1 0 51794 0 1 9891
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_0
timestamp 1666464484
transform 1 0 58128 0 1 20490
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_1
timestamp 1666464484
transform 1 0 58128 0 1 20146
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_2
timestamp 1666464484
transform 1 0 26187 0 1 19267
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_3
timestamp 1666464484
transform 1 0 26530 0 1 26206
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_4
timestamp 1666464484
transform 1 0 26545 0 1 19612
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_5
timestamp 1666464484
transform 1 0 27004 0 1 20490
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_6
timestamp 1666464484
transform 1 0 27004 0 1 20146
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_7
timestamp 1666464484
transform 1 0 24137 0 1 23593
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_8
timestamp 1666464484
transform 1 0 24149 0 1 17237
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_9
timestamp 1666464484
transform 1 0 24496 0 1 23915
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_10
timestamp 1666464484
transform 1 0 24509 0 1 17576
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_11
timestamp 1666464484
transform 1 0 24824 0 1 24236
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_12
timestamp 1666464484
transform 1 0 24837 0 1 17897
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_13
timestamp 1666464484
transform 1 0 25161 0 1 24557
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_14
timestamp 1666464484
transform 1 0 25174 0 1 18270
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_15
timestamp 1666464484
transform 1 0 25501 0 1 25248
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_16
timestamp 1666464484
transform 1 0 25514 0 1 18604
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_17
timestamp 1666464484
transform 1 0 25836 0 1 25567
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_18
timestamp 1666464484
transform 1 0 25851 0 1 18947
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_19
timestamp 1666464484
transform 1 0 26172 0 1 25887
box 0 0 1 1
use M3_M2431059054872_128x8m81  M3_M2431059054872_128x8m81_20
timestamp 1666464484
transform 1 0 41955 0 1 50533
box 0 0 1 1
use M3_M2431059054874_128x8m81  M3_M2431059054874_128x8m81_0
timestamp 1666464484
transform 1 0 43880 0 1 3016
box 0 0 1 1
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_0
timestamp 1666464484
transform 1 0 25674 0 1 51420
box -286 -162 286 162
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_1
timestamp 1666464484
transform 1 0 25674 0 1 31096
box -286 -162 286 162
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_2
timestamp 1666464484
transform 1 0 25674 0 1 30641
box -286 -162 286 162
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_3
timestamp 1666464484
transform 1 0 59149 0 1 31146
box -286 -162 286 162
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_4
timestamp 1666464484
transform 1 0 59149 0 1 30701
box -286 -162 286 162
use M3_M2431059054876_128x8m81  M3_M2431059054876_128x8m81_5
timestamp 1666464484
transform 1 0 59152 0 1 51420
box -286 -162 286 162
use M3_M2431059054878_128x8m81  M3_M2431059054878_128x8m81_0
timestamp 1666464484
transform 1 0 25660 0 1 34937
box -286 -348 286 348
use M3_M2431059054878_128x8m81  M3_M2431059054878_128x8m81_1
timestamp 1666464484
transform 1 0 59149 0 1 34906
box -286 -348 286 348
use M3_M2431059054879_128x8m81  M3_M2431059054879_128x8m81_0
timestamp 1666464484
transform 1 0 49313 0 1 1737
box -162 -472 162 472
use M3_M24310590548710_128x8m81  M3_M24310590548710_128x8m81_0
timestamp 1666464484
transform 1 0 48823 0 1 2670
box -162 -162 162 162
use M3_M24310590548714_128x8m81  M3_M24310590548714_128x8m81_0
timestamp 1666464484
transform 1 0 59135 0 1 27428
box -286 -906 286 906
use M3_M24310590548714_128x8m81  M3_M24310590548714_128x8m81_1
timestamp 1666464484
transform 1 0 25680 0 1 27367
box -286 -906 286 906
use M3_M24310590548718_128x8m81  M3_M24310590548718_128x8m81_0
timestamp 1666464484
transform 1 0 27590 0 1 34937
box -162 -348 162 348
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_0
timestamp 1666464484
transform 1 0 57495 0 1 22479
box -142 -454 142 454
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_1
timestamp 1666464484
transform 1 0 58126 0 1 23631
box -142 -454 142 454
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_2
timestamp 1666464484
transform 1 0 26990 0 1 23631
box -142 -454 142 454
use M3_M24310590548720_128x8m81  M3_M24310590548720_128x8m81_3
timestamp 1666464484
transform 1 0 27607 0 1 22492
box -142 -454 142 454
use control_512x8_128x8m81  control_512x8_128x8m81_0
timestamp 1666464484
transform 1 0 27533 0 1 4711
box -3624 -1833 31790 30125
use lcol4_128_128x8m81  lcol4_128_128x8m81_0
timestamp 1666464484
transform 1 0 2921 0 1 5019
box -1235 -3416 22810 46507
use m2m3_128x8m81  m2m3_128x8m81_0
timestamp 1666464484
transform 1 0 58611 0 1 17122
box 0 0 3541 9202
use power_a_128x8m81  power_a_128x8m81_0
timestamp 1666464484
transform -1 0 80818 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_1
timestamp 1666464484
transform 1 0 51233 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_2
timestamp 1666464484
transform 1 0 64218 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_3
timestamp 1666464484
transform 1 0 52478 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_4
timestamp 1666464484
transform 1 0 75018 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_5
timestamp 1666464484
transform 1 0 46033 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_6
timestamp 1666464484
transform 1 0 43633 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_7
timestamp 1666464484
transform -1 0 70018 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_8
timestamp 1666464484
transform -1 0 10442 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_9
timestamp 1666464484
transform -1 0 32324 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_10
timestamp 1666464484
transform -1 0 21242 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_11
timestamp 1666464484
transform -1 0 34022 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_12
timestamp 1666464484
transform 1 0 41233 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_13
timestamp 1666464484
transform 1 0 34831 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_14
timestamp 1666464484
transform 1 0 15442 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_15
timestamp 1666464484
transform 1 0 38028 0 1 282
box 0 -282 1000 1000
use power_a_128x8m81  power_a_128x8m81_16
timestamp 1666464484
transform 1 0 4642 0 1 282
box 0 -282 1000 1000
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_0
timestamp 1666464484
transform 1 0 15448 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_1
timestamp 1666464484
transform 1 0 10048 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_2
timestamp 1666464484
transform 1 0 4648 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_3
timestamp 1666464484
transform 1 0 64224 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_4
timestamp 1666464484
transform 1 0 69624 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_5
timestamp 1666464484
transform 1 0 75024 0 1 51346
box -511 630 1714 2430
use power_route_01_a_128x8m81  power_route_01_a_128x8m81_6
timestamp 1666464484
transform 1 0 46824 0 1 51346
box -511 630 1714 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_0
timestamp 1666464484
transform -1 0 21142 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_1
timestamp 1666464484
transform -1 0 41719 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_2
timestamp 1666464484
transform -1 0 80718 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_3
timestamp 1666464484
transform -1 0 85155 0 1 51346
box -511 630 489 2430
use power_route_01_b_128x8m81  power_route_01_b_128x8m81_4
timestamp 1666464484
transform -1 0 45558 0 1 51346
box -511 630 489 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_0
timestamp 1666464484
transform -1 0 34095 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_1
timestamp 1666464484
transform -1 0 38662 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_2
timestamp 1666464484
transform -1 0 30987 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_3
timestamp 1666464484
transform -1 0 29591 0 1 51346
box 714 1822 1714 2430
use power_route_01_c_128x8m81  power_route_01_c_128x8m81_4
timestamp 1666464484
transform -1 0 44144 0 1 51346
box 714 1822 1714 2430
use power_route_128_128x8m81  power_route_128_128x8m81_0
timestamp 1666464484
transform 1 0 -1921 0 1 -2063
box 1921 2345 88293 55839
use rcol4_128_128x8m81  rcol4_128_128x8m81_0
timestamp 1666464484
transform 1 0 60511 0 1 5019
box -1090 -3398 24602 46517
use xdec16_128_128x8m81  xdec16_128_128x8m81_0
timestamp 1666464484
transform 1 0 28677 0 1 36127
box -3364 -228 31133 15548
<< labels >>
flabel metal3 s 2626 53168 3626 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 50176 1706 50876 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 48376 1706 49076 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 4642 0 5642 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 5362 53168 6362 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 46576 1706 47276 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 44776 1706 45476 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 8026 53168 9026 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 42976 1706 43676 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 41176 1706 41876 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 39376 1706 40076 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 37576 1706 38276 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 9442 0 10442 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 35776 1706 36476 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 8152 3011 9515 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 10762 53168 11762 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 8153 24250 9515 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 13426 53168 14426 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 15442 0 16442 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 16162 53168 17162 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 28178 7084 28729 9516 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 24047 8154 28729 9516 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29537 6744 34622 7652 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 18826 53168 19826 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 20242 0 21242 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 28178 7084 34622 7652 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 22258 53168 23258 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 25158 53168 26158 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 1401 51976 2401 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 4137 51976 5137 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 34536 27828 35326 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 6801 51976 7801 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 6921 26434 8163 28416 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 17721 26434 18963 28416 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 26435 26070 28416 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 9537 51976 10537 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 26435 27828 26890 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 12201 51976 13201 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 14937 51976 15937 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 10176 3011 11493 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 2249 10174 24250 11491 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 17601 51976 18601 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 20653 51976 21653 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 2229 10175 24250 11491 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 24047 10176 27828 11493 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 27877 53168 28877 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29273 53168 30273 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 23483 51976 24483 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 31324 0 32324 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26572 51976 27572 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 32381 53168 33381 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 30710 51976 31710 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 35415 51976 36415 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 33022 0 34022 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 38585 51976 39585 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 34024 53168 35024 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 34831 0 35831 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 41230 51976 42230 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 45069 51976 46069 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 36948 53168 37948 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 38028 0 39028 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 39882 53168 40882 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 46313 51976 47313 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 41233 0 42233 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 42430 53168 43430 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 48901 51976 49901 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 52569 51976 53569 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 54262 51976 55262 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 43633 0 44633 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 43713 53168 44713 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 57547 51976 58547 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 60977 51976 61977 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 46033 0 47033 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 47538 53168 48538 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 63713 51976 64713 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50465 53168 51465 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 66377 51976 67377 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 51233 0 52233 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 69113 51976 70113 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 71777 51976 72777 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 52478 0 53478 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 55990 53168 56990 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 74513 51976 75513 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 77177 51976 78177 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 80229 51976 81229 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 83059 51976 84059 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 51976 85666 53776 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51976 86372 52976 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 50176 86372 50876 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 53168 59791 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 62202 53168 63202 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 64218 0 65218 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 48376 86372 49076 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 64938 53168 65938 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 67602 53168 68602 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 46576 86372 47276 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 69018 0 70018 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 70338 53168 71338 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 44776 86372 45476 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 42976 86372 43676 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 73002 53168 74002 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 75018 0 76018 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 75738 53168 76738 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 41176 86372 41876 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 78402 53168 79402 53776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 39376 86372 40076 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 79818 0 80818 932 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 37576 86372 38276 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 81834 53168 82834 53776 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 84666 35776 86372 36476 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 29430 1706 34125 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 2095 32315 2188 34126 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51076 1014 51776 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 32315 3011 34125 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 32316 25085 34125 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51226 27779 51626 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 32318 27214 34124 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 26772 31486 58351 32199 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30402 51326 54622 51528 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26772 27382 58351 30105 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 31486 58351 34124 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61853 32315 72383 34125 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 32315 86372 34124 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 51327 86372 51528 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 29430 86372 29714 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 29430 86372 34125 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 51258 59517 51591 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 72653 32315 86372 34125 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 58791 51276 86372 51576 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 22938 1706 23938 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 85358 51076 86372 51776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 22938 27214 23380 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 49276 1014 49976 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26770 23370 58348 24278 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 22937 83763 23380 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57908 22938 86372 23380 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 22938 86372 23938 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 18016 24250 20739 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 49476 27272 49776 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29513 19969 55645 21625 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 49526 54622 49728 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 49526 86372 49726 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 49476 86372 49776 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 85358 49276 86372 49976 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 29521 19969 55645 21707 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 44432 19969 55645 21708 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61825 18015 83763 20739 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61807 18016 86372 20739 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 19969 86372 20739 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 47476 1014 48176 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 47676 27272 47976 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 12036 1706 14178 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 23821 12046 34761 12847 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 13461 27214 14178 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 12036 24250 12846 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 24047 12046 27214 14179 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 47726 54622 47928 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 24047 12046 34761 12934 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 34741 9972 41516 12574 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29478 10756 41516 12574 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 29478 11697 58351 12574 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 47726 86372 47926 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 47676 86372 47976 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 85358 47476 86372 48176 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 45676 1014 46376 0 FreeSans 2000 180 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 26772 11844 58351 12574 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 12035 58421 13866 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 59826 12035 60026 14017 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 13461 86372 13866 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61807 13461 72429 14178 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61773 13461 86372 14177 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 83169 12035 84221 12847 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 45876 27272 46176 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 83169 13461 84221 14179 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 50228 12036 86372 12846 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 26772 12035 84999 12574 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 84666 12036 86372 14178 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 72607 13461 86372 14178 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61802 8153 86372 9514 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 57909 8154 62278 9516 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 61825 8152 86372 9514 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 30403 45926 54622 46128 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 83361 8152 86372 9515 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 45926 86372 46126 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 59421 45876 86372 46176 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 4060 1712 5629 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 85358 45676 86372 46376 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 5173 3011 5629 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 43876 1014 44576 0 FreeSans 2000 0 0 0 VSS
port 28 nsew ground bidirectional
flabel metal3 s 0 5174 24250 5629 0 FreeSans 2000 0 0 0 VDD
port 27 nsew power bidirectional
flabel metal3 s 0 4060 24341 4515 0 FreeSans 2000 180 0 0 VDD
port 27 nsew power bidirectional
rlabel metal2 s 27936 0 28160 200 4 CLK
port 9 nsew signal input
rlabel metal2 s 1864 0 2088 200 4 D[0]
port 17 nsew signal input
rlabel metal2 s 30859 0 31083 200 4 A[2]
port 5 nsew signal input
rlabel metal2 s 32552 0 32776 200 4 A[1]
port 6 nsew signal input
rlabel metal2 s 34243 0 34467 200 4 A[0]
port 7 nsew signal input
rlabel metal2 s 14127 0 14351 200 4 Q[2]
port 24 nsew signal output
rlabel metal2 s 22279 0 22503 200 4 Q[3]
port 23 nsew signal output
rlabel metal2 s 50342 0 50566 200 4 CEN
port 8 nsew signal input
rlabel metal2 s 54417 0 54641 200 4 A[5]
port 2 nsew signal input
rlabel metal2 s 53772 0 53996 200 4 A[6]
port 1 nsew signal input
rlabel metal2 s 55164 0 55388 200 4 A[4]
port 3 nsew signal input
rlabel metal2 s 23404 0 23628 200 4 WEN[3]
port 33 nsew signal input
rlabel metal2 s 83372 0 83596 200 4 D[7]
port 10 nsew signal input
rlabel metal2 s 81855 0 82079 200 4 Q[7]
port 19 nsew signal output
rlabel metal2 s 23795 0 24019 200 4 D[3]
port 14 nsew signal input
rlabel metal2 s 12206 0 12430 200 4 D[1]
port 16 nsew signal input
rlabel metal2 s 13454 0 13678 200 4 D[2]
port 15 nsew signal input
rlabel metal2 s 56265 0 56489 200 4 A[3]
port 4 nsew signal input
rlabel metal2 s 11533 0 11757 200 4 Q[1]
port 25 nsew signal output
rlabel metal2 s 73703 0 73927 200 4 Q[6]
port 20 nsew signal output
rlabel metal2 s 71782 0 72006 200 4 D[5]
port 12 nsew signal input
rlabel metal2 s 62958 0 63182 200 4 Q[4]
port 22 nsew signal output
rlabel metal2 s 72180 0 72404 200 4 WEN[5]
port 31 nsew signal input
rlabel metal2 s 13054 0 13278 200 4 WEN[2]
port 34 nsew signal input
rlabel metal2 s 12604 0 12828 200 4 WEN[1]
port 35 nsew signal input
rlabel metal2 s 62115 0 62339 200 4 WEN[4]
port 32 nsew signal input
rlabel metal2 s 82695 0 82919 200 4 WEN[7]
port 29 nsew signal input
rlabel metal2 s 72630 0 72854 200 4 WEN[6]
port 30 nsew signal input
rlabel metal2 s 61447 0 61671 200 4 D[4]
port 13 nsew signal input
rlabel metal2 s 73030 0 73254 200 4 D[6]
port 11 nsew signal input
rlabel metal2 s 71109 0 71333 200 4 Q[5]
port 21 nsew signal output
rlabel metal2 s 3380 0 3604 200 4 Q[0]
port 26 nsew signal output
rlabel metal2 s 40588 0 40812 200 4 GWEN
port 18 nsew signal input
rlabel metal2 s 2539 0 2763 200 4 WEN[0]
port 36 nsew signal input
flabel space 0 200 0 200 3 FreeSans 2000 0 0 0 & Metric 1.00
flabel space 0 600 0 600 3 FreeSans 2000 0 0 0 & Version 2015q2v1
flabel space 0 1000 0 1000 3 FreeSans 2000 0 0 0 & Product GF018_5VGreen_SRAM_1P_128x8M8WM1
flabel metal3 0 1400 0 1400 3 FreeSans 2000 0 0 0 & Vendor GLOBALFOUNDRIES
rlabel metal3 s 23687 5175 27214 5630 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23909 4166 62429 4619 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 4164 59323 4515 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 4166 62429 4621 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57909 5175 62429 5630 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61788 4060 86372 4515 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 83361 5173 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 61802 5174 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84660 4060 86372 5629 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 706 0 1706 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 2039 0 3039 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 3442 0 4442 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 5842 0 6842 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 7042 0 8042 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 8242 0 9242 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 10642 0 11642 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 12443 0 13443 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 14242 0 15242 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 16642 0 17642 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 17842 0 18842 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 19042 0 20042 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 21910 0 22910 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 23110 0 24110 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 24410 0 25410 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 25710 0 26710 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 27010 0 28010 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 28310 0 29310 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 29610 0 30610 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 36031 0 37031 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 39228 0 40228 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 42433 0 43433 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 44833 0 45833 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 47233 0 48233 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 48566 0 49566 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 49876 0 50876 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 54458 0 55458 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 55758 0 56758 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 57058 0 58058 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 58358 0 59358 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 59658 0 60658 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 60958 0 61958 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 62295 0 63295 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 65418 0 66418 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 66618 0 67618 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 67818 0 68818 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 70218 0 71218 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 72017 0 73017 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 73818 0 74818 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 76218 0 77218 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 77418 0 78418 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 78618 0 79618 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 81018 0 82018 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 82419 0 83419 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 84666 0 85666 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 1232 86372 2232 1 VDD
port 27 nsew power bidirectional
rlabel metal3 s 0 44076 27272 44376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 44126 54622 44328 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 44126 86372 44326 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 44076 86372 44376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 43876 86372 44576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42076 1014 42776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42276 27272 42576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 42326 54622 42528 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 42326 86372 42526 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 42276 86372 42576 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 42076 86372 42776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40276 1014 40976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40476 27272 40776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 40526 54622 40728 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 40526 86372 40726 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 40476 86372 40776 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 40276 86372 40976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38476 1014 39176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38676 27272 38976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 38726 54622 38928 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 38726 86372 38926 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 38676 86372 38976 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 38476 86372 39176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36676 1014 37376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36876 27272 37176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 30403 36926 54622 37128 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 36926 86372 37126 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 59421 36876 86372 37176 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 36676 86372 37376 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57369 34536 86372 35326 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 26435 86372 26890 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 66497 26434 67739 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 77297 26434 78539 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 58785 26435 86372 28416 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21282 1014 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24036 21826 27826 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 21827 27826 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 21826 27826 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 57677 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 22291 57677 23199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21826 83763 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 21282 86372 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 56078 21827 86372 22282 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 23678 17730 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14328 24250 16597 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 24111 14329 27828 16598 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29478 13243 45977 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27387 13245 45977 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14491 47683 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41493 13078 49775 13760 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14936 51760 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 14966 55645 15015 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46982 14968 86372 16784 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 14327 83763 16784 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61807 14328 86372 17730 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42261 10740 57736 11527 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 10176 86372 11491 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10173 84482 11493 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61805 10175 84482 11491 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 10176 86372 11493 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 1014 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 3011 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 6982 3011 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2249 6980 24250 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 2226 6981 24250 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23625 6982 27828 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23687 6177 41397 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 5665 34622 6573 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 5766 34622 6198 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29458 6177 41397 6573 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6177 41397 8582 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 29513 7900 41397 8582 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 34860 6592 55482 7392 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41857 9165 51430 10420 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5605 55482 9502 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 57736 8888 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57295 6982 86372 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 62429 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 6984 62747 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 50922 5766 86372 6198 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61825 6980 84787 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 61802 6981 84787 7595 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 5766 86372 6199 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 5766 86372 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 83361 6982 86372 7596 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 1000 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3420 3011 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 3421 24341 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 27438 3524 27778 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 28764 3524 28894 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 41774 3524 41904 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 42299 3524 42429 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 46873 3524 47003 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47321 3524 47451 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 47769 3524 47899 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 48217 3524 48347 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 23909 3524 61215 3875 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 57345 3524 61215 3876 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 0 2502 86372 2854 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 60886 3420 86372 3772 1 VSS
port 28 nsew ground bidirectional
rlabel metal3 s 85358 2502 86372 3772 1 VSS
port 28 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 86372 53776
string GDS_END 2348210
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2298636
string LEFclass BLOCK
string LEFsymmetry X Y R90
string path 307.290 11.160 307.290 0.000 
<< end >>
