magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 2344 664
<< mvpmos >>
rect 0 0 120 544
rect 224 0 344 544
rect 448 0 568 544
rect 672 0 792 544
rect 896 0 1016 544
rect 1120 0 1240 544
rect 1344 0 1464 544
rect 1568 0 1688 544
rect 1792 0 1912 544
rect 2016 0 2136 544
<< mvpdiff >>
rect -88 531 0 544
rect -88 485 -75 531
rect -29 485 0 531
rect -88 413 0 485
rect -88 367 -75 413
rect -29 367 0 413
rect -88 295 0 367
rect -88 249 -75 295
rect -29 249 0 295
rect -88 177 0 249
rect -88 131 -75 177
rect -29 131 0 177
rect -88 59 0 131
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 531 224 544
rect 120 485 149 531
rect 195 485 224 531
rect 120 413 224 485
rect 120 367 149 413
rect 195 367 224 413
rect 120 295 224 367
rect 120 249 149 295
rect 195 249 224 295
rect 120 177 224 249
rect 120 131 149 177
rect 195 131 224 177
rect 120 59 224 131
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 531 448 544
rect 344 485 373 531
rect 419 485 448 531
rect 344 413 448 485
rect 344 367 373 413
rect 419 367 448 413
rect 344 295 448 367
rect 344 249 373 295
rect 419 249 448 295
rect 344 177 448 249
rect 344 131 373 177
rect 419 131 448 177
rect 344 59 448 131
rect 344 13 373 59
rect 419 13 448 59
rect 344 0 448 13
rect 568 531 672 544
rect 568 485 597 531
rect 643 485 672 531
rect 568 413 672 485
rect 568 367 597 413
rect 643 367 672 413
rect 568 295 672 367
rect 568 249 597 295
rect 643 249 672 295
rect 568 177 672 249
rect 568 131 597 177
rect 643 131 672 177
rect 568 59 672 131
rect 568 13 597 59
rect 643 13 672 59
rect 568 0 672 13
rect 792 531 896 544
rect 792 485 821 531
rect 867 485 896 531
rect 792 413 896 485
rect 792 367 821 413
rect 867 367 896 413
rect 792 295 896 367
rect 792 249 821 295
rect 867 249 896 295
rect 792 177 896 249
rect 792 131 821 177
rect 867 131 896 177
rect 792 59 896 131
rect 792 13 821 59
rect 867 13 896 59
rect 792 0 896 13
rect 1016 531 1120 544
rect 1016 485 1045 531
rect 1091 485 1120 531
rect 1016 413 1120 485
rect 1016 367 1045 413
rect 1091 367 1120 413
rect 1016 295 1120 367
rect 1016 249 1045 295
rect 1091 249 1120 295
rect 1016 177 1120 249
rect 1016 131 1045 177
rect 1091 131 1120 177
rect 1016 59 1120 131
rect 1016 13 1045 59
rect 1091 13 1120 59
rect 1016 0 1120 13
rect 1240 531 1344 544
rect 1240 485 1269 531
rect 1315 485 1344 531
rect 1240 413 1344 485
rect 1240 367 1269 413
rect 1315 367 1344 413
rect 1240 295 1344 367
rect 1240 249 1269 295
rect 1315 249 1344 295
rect 1240 177 1344 249
rect 1240 131 1269 177
rect 1315 131 1344 177
rect 1240 59 1344 131
rect 1240 13 1269 59
rect 1315 13 1344 59
rect 1240 0 1344 13
rect 1464 531 1568 544
rect 1464 485 1493 531
rect 1539 485 1568 531
rect 1464 413 1568 485
rect 1464 367 1493 413
rect 1539 367 1568 413
rect 1464 295 1568 367
rect 1464 249 1493 295
rect 1539 249 1568 295
rect 1464 177 1568 249
rect 1464 131 1493 177
rect 1539 131 1568 177
rect 1464 59 1568 131
rect 1464 13 1493 59
rect 1539 13 1568 59
rect 1464 0 1568 13
rect 1688 531 1792 544
rect 1688 485 1717 531
rect 1763 485 1792 531
rect 1688 413 1792 485
rect 1688 367 1717 413
rect 1763 367 1792 413
rect 1688 295 1792 367
rect 1688 249 1717 295
rect 1763 249 1792 295
rect 1688 177 1792 249
rect 1688 131 1717 177
rect 1763 131 1792 177
rect 1688 59 1792 131
rect 1688 13 1717 59
rect 1763 13 1792 59
rect 1688 0 1792 13
rect 1912 531 2016 544
rect 1912 485 1941 531
rect 1987 485 2016 531
rect 1912 413 2016 485
rect 1912 367 1941 413
rect 1987 367 2016 413
rect 1912 295 2016 367
rect 1912 249 1941 295
rect 1987 249 2016 295
rect 1912 177 2016 249
rect 1912 131 1941 177
rect 1987 131 2016 177
rect 1912 59 2016 131
rect 1912 13 1941 59
rect 1987 13 2016 59
rect 1912 0 2016 13
rect 2136 531 2224 544
rect 2136 485 2165 531
rect 2211 485 2224 531
rect 2136 413 2224 485
rect 2136 367 2165 413
rect 2211 367 2224 413
rect 2136 295 2224 367
rect 2136 249 2165 295
rect 2211 249 2224 295
rect 2136 177 2224 249
rect 2136 131 2165 177
rect 2211 131 2224 177
rect 2136 59 2224 131
rect 2136 13 2165 59
rect 2211 13 2224 59
rect 2136 0 2224 13
<< mvpdiffc >>
rect -75 485 -29 531
rect -75 367 -29 413
rect -75 249 -29 295
rect -75 131 -29 177
rect -75 13 -29 59
rect 149 485 195 531
rect 149 367 195 413
rect 149 249 195 295
rect 149 131 195 177
rect 149 13 195 59
rect 373 485 419 531
rect 373 367 419 413
rect 373 249 419 295
rect 373 131 419 177
rect 373 13 419 59
rect 597 485 643 531
rect 597 367 643 413
rect 597 249 643 295
rect 597 131 643 177
rect 597 13 643 59
rect 821 485 867 531
rect 821 367 867 413
rect 821 249 867 295
rect 821 131 867 177
rect 821 13 867 59
rect 1045 485 1091 531
rect 1045 367 1091 413
rect 1045 249 1091 295
rect 1045 131 1091 177
rect 1045 13 1091 59
rect 1269 485 1315 531
rect 1269 367 1315 413
rect 1269 249 1315 295
rect 1269 131 1315 177
rect 1269 13 1315 59
rect 1493 485 1539 531
rect 1493 367 1539 413
rect 1493 249 1539 295
rect 1493 131 1539 177
rect 1493 13 1539 59
rect 1717 485 1763 531
rect 1717 367 1763 413
rect 1717 249 1763 295
rect 1717 131 1763 177
rect 1717 13 1763 59
rect 1941 485 1987 531
rect 1941 367 1987 413
rect 1941 249 1987 295
rect 1941 131 1987 177
rect 1941 13 1987 59
rect 2165 485 2211 531
rect 2165 367 2211 413
rect 2165 249 2211 295
rect 2165 131 2211 177
rect 2165 13 2211 59
<< polysilicon >>
rect 0 544 120 588
rect 224 544 344 588
rect 448 544 568 588
rect 672 544 792 588
rect 896 544 1016 588
rect 1120 544 1240 588
rect 1344 544 1464 588
rect 1568 544 1688 588
rect 1792 544 1912 588
rect 2016 544 2136 588
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
<< metal1 >>
rect -75 531 -29 544
rect -75 413 -29 485
rect -75 295 -29 367
rect -75 177 -29 249
rect -75 59 -29 131
rect -75 0 -29 13
rect 149 531 195 544
rect 149 413 195 485
rect 149 295 195 367
rect 149 177 195 249
rect 149 59 195 131
rect 149 0 195 13
rect 373 531 419 544
rect 373 413 419 485
rect 373 295 419 367
rect 373 177 419 249
rect 373 59 419 131
rect 373 0 419 13
rect 597 531 643 544
rect 597 413 643 485
rect 597 295 643 367
rect 597 177 643 249
rect 597 59 643 131
rect 597 0 643 13
rect 821 531 867 544
rect 821 413 867 485
rect 821 295 867 367
rect 821 177 867 249
rect 821 59 867 131
rect 821 0 867 13
rect 1045 531 1091 544
rect 1045 413 1091 485
rect 1045 295 1091 367
rect 1045 177 1091 249
rect 1045 59 1091 131
rect 1045 0 1091 13
rect 1269 531 1315 544
rect 1269 413 1315 485
rect 1269 295 1315 367
rect 1269 177 1315 249
rect 1269 59 1315 131
rect 1269 0 1315 13
rect 1493 531 1539 544
rect 1493 413 1539 485
rect 1493 295 1539 367
rect 1493 177 1539 249
rect 1493 59 1539 131
rect 1493 0 1539 13
rect 1717 531 1763 544
rect 1717 413 1763 485
rect 1717 295 1763 367
rect 1717 177 1763 249
rect 1717 59 1763 131
rect 1717 0 1763 13
rect 1941 531 1987 544
rect 1941 413 1987 485
rect 1941 295 1987 367
rect 1941 177 1987 249
rect 1941 59 1987 131
rect 1941 0 1987 13
rect 2165 531 2211 544
rect 2165 413 2211 485
rect 2165 295 2211 367
rect 2165 177 2211 249
rect 2165 59 2211 131
rect 2165 0 2211 13
<< labels >>
flabel metal1 s -52 272 -52 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 2188 272 2188 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 272 172 272 0 FreeSans 400 0 0 0 D
flabel metal1 s 396 272 396 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 620 272 620 272 0 FreeSans 400 0 0 0 D
flabel metal1 s 844 272 844 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 1068 272 1068 272 0 FreeSans 400 0 0 0 D
flabel metal1 s 1292 272 1292 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 1516 272 1516 272 0 FreeSans 400 0 0 0 D
flabel metal1 s 1740 272 1740 272 0 FreeSans 400 0 0 0 S
flabel metal1 s 1964 272 1964 272 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 45998
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 38080
<< end >>
