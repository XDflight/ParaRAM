magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -1734 23 1734 42
rect -1734 -23 -1715 23
rect 1715 -23 1734 23
rect -1734 -42 1734 -23
<< psubdiffcont >>
rect -1715 -23 1715 23
<< metal1 >>
rect -1726 23 1726 34
rect -1726 -23 -1715 23
rect 1715 -23 1726 23
rect -1726 -34 1726 -23
<< properties >>
string GDS_END 1804474
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1801910
<< end >>
