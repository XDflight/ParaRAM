magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 11494 14188 11623 14228
rect 11494 14136 11532 14188
rect 11584 14136 11623 14188
rect 11494 14109 11623 14136
rect 11494 14096 11622 14109
rect 12627 13957 12756 13997
rect 12627 13905 12665 13957
rect 12717 13905 12756 13957
rect 12627 13878 12756 13905
rect 12627 13865 12755 13878
rect 15156 13848 15285 13888
rect 15156 13796 15194 13848
rect 15246 13796 15285 13848
rect 15156 13769 15285 13796
rect 15156 13756 15284 13769
rect 15534 13204 15663 13244
rect 15534 13152 15572 13204
rect 15624 13152 15663 13204
rect 12627 13095 12756 13135
rect 15534 13125 15663 13152
rect 15534 13112 15662 13125
rect 12627 13043 12665 13095
rect 12717 13043 12756 13095
rect 12627 13016 12756 13043
rect 12627 13003 12755 13016
rect 11494 12864 11623 12904
rect 11494 12812 11532 12864
rect 11584 12812 11623 12864
rect 11494 12785 11623 12812
rect 11494 12772 11622 12785
rect 11494 12388 11623 12428
rect 11494 12336 11532 12388
rect 11584 12336 11623 12388
rect 11494 12309 11623 12336
rect 11494 12296 11622 12309
rect 12627 12157 12756 12197
rect 12627 12105 12665 12157
rect 12717 12105 12756 12157
rect 12627 12078 12756 12105
rect 12627 12065 12755 12078
rect 15912 12048 16041 12088
rect 15912 11996 15950 12048
rect 16002 11996 16041 12048
rect 15912 11969 16041 11996
rect 15912 11956 16040 11969
rect 16290 11404 16419 11444
rect 16290 11352 16328 11404
rect 16380 11352 16419 11404
rect 12627 11295 12756 11335
rect 16290 11325 16419 11352
rect 16290 11312 16418 11325
rect 12627 11243 12665 11295
rect 12717 11243 12756 11295
rect 12627 11216 12756 11243
rect 12627 11203 12755 11216
rect 11494 11064 11623 11104
rect 11494 11012 11532 11064
rect 11584 11012 11623 11064
rect 11494 10985 11623 11012
rect 11494 10972 11622 10985
rect 11494 10588 11623 10628
rect 11494 10536 11532 10588
rect 11584 10536 11623 10588
rect 11494 10509 11623 10536
rect 11494 10496 11622 10509
rect 12627 10357 12756 10397
rect 12627 10305 12665 10357
rect 12717 10305 12756 10357
rect 12627 10278 12756 10305
rect 12627 10265 12755 10278
rect 16667 10248 16796 10288
rect 16667 10196 16705 10248
rect 16757 10196 16796 10248
rect 16667 10169 16796 10196
rect 16667 10156 16795 10169
rect 17045 9604 17174 9644
rect 17045 9552 17083 9604
rect 17135 9552 17174 9604
rect 12627 9495 12756 9535
rect 17045 9525 17174 9552
rect 17045 9512 17173 9525
rect 12627 9443 12665 9495
rect 12717 9443 12756 9495
rect 12627 9416 12756 9443
rect 12627 9403 12755 9416
rect 11494 9264 11623 9304
rect 11494 9212 11532 9264
rect 11584 9212 11623 9264
rect 11494 9185 11623 9212
rect 11494 9172 11622 9185
rect 11494 8788 11623 8828
rect 11494 8736 11532 8788
rect 11584 8736 11623 8788
rect 11494 8709 11623 8736
rect 11494 8696 11622 8709
rect 12627 8557 12756 8597
rect 12627 8505 12665 8557
rect 12717 8505 12756 8557
rect 12627 8478 12756 8505
rect 12627 8465 12755 8478
rect 17423 8448 17552 8488
rect 17423 8396 17461 8448
rect 17513 8396 17552 8448
rect 17423 8369 17552 8396
rect 17423 8356 17551 8369
rect 17800 7804 17929 7844
rect 17800 7752 17838 7804
rect 17890 7752 17929 7804
rect 12627 7695 12756 7735
rect 17800 7725 17929 7752
rect 17800 7712 17928 7725
rect 12627 7643 12665 7695
rect 12717 7643 12756 7695
rect 12627 7616 12756 7643
rect 12627 7603 12755 7616
rect 11494 7464 11623 7504
rect 11494 7412 11532 7464
rect 11584 7412 11623 7464
rect 11494 7385 11623 7412
rect 11494 7372 11622 7385
rect 11494 6988 11623 7028
rect 11494 6936 11532 6988
rect 11584 6936 11623 6988
rect 11494 6909 11623 6936
rect 11494 6896 11622 6909
rect 13004 6757 13133 6797
rect 13004 6705 13042 6757
rect 13094 6705 13133 6757
rect 13004 6678 13133 6705
rect 13004 6665 13132 6678
rect 15156 6648 15285 6688
rect 15156 6596 15194 6648
rect 15246 6596 15285 6648
rect 15156 6569 15285 6596
rect 15156 6556 15284 6569
rect 15534 6004 15663 6044
rect 15534 5952 15572 6004
rect 15624 5952 15663 6004
rect 13004 5895 13133 5935
rect 15534 5925 15663 5952
rect 15534 5912 15662 5925
rect 13004 5843 13042 5895
rect 13094 5843 13133 5895
rect 13004 5816 13133 5843
rect 13004 5803 13132 5816
rect 11494 5664 11623 5704
rect 11494 5612 11532 5664
rect 11584 5612 11623 5664
rect 11494 5585 11623 5612
rect 11494 5572 11622 5585
rect 11494 5188 11623 5228
rect 11494 5136 11532 5188
rect 11584 5136 11623 5188
rect 11494 5109 11623 5136
rect 11494 5096 11622 5109
rect 13004 4957 13133 4997
rect 13004 4905 13042 4957
rect 13094 4905 13133 4957
rect 13004 4878 13133 4905
rect 13004 4865 13132 4878
rect 15912 4848 16041 4888
rect 15912 4796 15950 4848
rect 16002 4796 16041 4848
rect 15912 4769 16041 4796
rect 15912 4756 16040 4769
rect 16290 4204 16419 4244
rect 16290 4152 16328 4204
rect 16380 4152 16419 4204
rect 13004 4095 13133 4135
rect 16290 4125 16419 4152
rect 16290 4112 16418 4125
rect 13004 4043 13042 4095
rect 13094 4043 13133 4095
rect 13004 4016 13133 4043
rect 13004 4003 13132 4016
rect 11494 3864 11623 3904
rect 11494 3812 11532 3864
rect 11584 3812 11623 3864
rect 11494 3785 11623 3812
rect 11494 3772 11622 3785
rect 11494 3388 11623 3428
rect 11494 3336 11532 3388
rect 11584 3336 11623 3388
rect 11494 3309 11623 3336
rect 11494 3296 11622 3309
rect 13004 3157 13133 3197
rect 13004 3105 13042 3157
rect 13094 3105 13133 3157
rect 13004 3078 13133 3105
rect 13004 3065 13132 3078
rect 16667 3048 16796 3088
rect 16667 2996 16705 3048
rect 16757 2996 16796 3048
rect 16667 2969 16796 2996
rect 16667 2956 16795 2969
rect 17045 2404 17174 2444
rect 17045 2352 17083 2404
rect 17135 2352 17174 2404
rect 13004 2295 13133 2335
rect 17045 2325 17174 2352
rect 17045 2312 17173 2325
rect 13004 2243 13042 2295
rect 13094 2243 13133 2295
rect 13004 2216 13133 2243
rect 13004 2203 13132 2216
rect 11494 2064 11623 2104
rect 11494 2012 11532 2064
rect 11584 2012 11623 2064
rect 11494 1985 11623 2012
rect 11494 1972 11622 1985
rect 11494 1588 11623 1628
rect 11494 1536 11532 1588
rect 11584 1536 11623 1588
rect 11494 1509 11623 1536
rect 11494 1496 11622 1509
rect 13004 1357 13133 1397
rect 13004 1305 13042 1357
rect 13094 1305 13133 1357
rect 13004 1278 13133 1305
rect 13004 1265 13132 1278
rect 17423 1248 17552 1288
rect 17423 1196 17461 1248
rect 17513 1196 17552 1248
rect 17423 1169 17552 1196
rect 17423 1156 17551 1169
rect 17800 604 17929 644
rect 17800 552 17838 604
rect 17890 552 17929 604
rect 13004 495 13133 535
rect 17800 525 17929 552
rect 17800 512 17928 525
rect 13004 443 13042 495
rect 13094 443 13133 495
rect 13004 416 13133 443
rect 13004 403 13132 416
rect 11494 264 11623 304
rect 11494 212 11532 264
rect 11584 212 11623 264
rect 11494 185 11623 212
rect 11494 172 11622 185
<< via1 >>
rect 11532 14136 11584 14188
rect 12665 13905 12717 13957
rect 15194 13796 15246 13848
rect 15572 13152 15624 13204
rect 12665 13043 12717 13095
rect 11532 12812 11584 12864
rect 11532 12336 11584 12388
rect 12665 12105 12717 12157
rect 15950 11996 16002 12048
rect 16328 11352 16380 11404
rect 12665 11243 12717 11295
rect 11532 11012 11584 11064
rect 11532 10536 11584 10588
rect 12665 10305 12717 10357
rect 16705 10196 16757 10248
rect 17083 9552 17135 9604
rect 12665 9443 12717 9495
rect 11532 9212 11584 9264
rect 11532 8736 11584 8788
rect 12665 8505 12717 8557
rect 17461 8396 17513 8448
rect 17838 7752 17890 7804
rect 12665 7643 12717 7695
rect 11532 7412 11584 7464
rect 11532 6936 11584 6988
rect 13042 6705 13094 6757
rect 15194 6596 15246 6648
rect 15572 5952 15624 6004
rect 13042 5843 13094 5895
rect 11532 5612 11584 5664
rect 11532 5136 11584 5188
rect 13042 4905 13094 4957
rect 15950 4796 16002 4848
rect 16328 4152 16380 4204
rect 13042 4043 13094 4095
rect 11532 3812 11584 3864
rect 11532 3336 11584 3388
rect 13042 3105 13094 3157
rect 16705 2996 16757 3048
rect 17083 2352 17135 2404
rect 13042 2243 13094 2295
rect 11532 2012 11584 2064
rect 11532 1536 11584 1588
rect 13042 1305 13094 1357
rect 17461 1196 17513 1248
rect 17838 552 17890 604
rect 13042 443 13094 495
rect 11532 212 11584 264
<< metal2 >>
rect 11494 14188 11622 14229
rect 11494 14136 11532 14188
rect 11584 14136 11622 14188
rect 11494 14095 11622 14136
rect 12627 13957 12755 13998
rect 12627 13905 12665 13957
rect 12717 13905 12755 13957
rect 12627 13864 12755 13905
rect 15156 13848 15284 13889
rect 15156 13796 15194 13848
rect 15246 13796 15284 13848
rect 15156 13755 15284 13796
rect 15534 13204 15662 13245
rect 15534 13152 15572 13204
rect 15624 13152 15662 13204
rect 12627 13095 12755 13136
rect 15534 13111 15662 13152
rect 12627 13043 12665 13095
rect 12717 13043 12755 13095
rect 12627 13002 12755 13043
rect 11494 12864 11622 12905
rect 11494 12812 11532 12864
rect 11584 12812 11622 12864
rect 11494 12771 11622 12812
rect 11494 12388 11622 12429
rect 11494 12336 11532 12388
rect 11584 12336 11622 12388
rect 11494 12295 11622 12336
rect 12627 12157 12755 12198
rect 12627 12105 12665 12157
rect 12717 12105 12755 12157
rect 12627 12064 12755 12105
rect 15912 12048 16040 12089
rect 15912 11996 15950 12048
rect 16002 11996 16040 12048
rect 15912 11955 16040 11996
rect 16290 11404 16418 11445
rect 16290 11352 16328 11404
rect 16380 11352 16418 11404
rect 12627 11295 12755 11336
rect 16290 11311 16418 11352
rect 12627 11243 12665 11295
rect 12717 11243 12755 11295
rect 12627 11202 12755 11243
rect 11494 11064 11622 11105
rect 11494 11012 11532 11064
rect 11584 11012 11622 11064
rect 11494 10971 11622 11012
rect 11494 10588 11622 10629
rect 11494 10536 11532 10588
rect 11584 10536 11622 10588
rect 11494 10495 11622 10536
rect 12627 10357 12755 10398
rect 12627 10305 12665 10357
rect 12717 10305 12755 10357
rect 12627 10264 12755 10305
rect 16667 10248 16795 10289
rect 16667 10196 16705 10248
rect 16757 10196 16795 10248
rect 16667 10155 16795 10196
rect 17045 9604 17173 9645
rect 17045 9552 17083 9604
rect 17135 9552 17173 9604
rect 12627 9495 12755 9536
rect 17045 9511 17173 9552
rect 12627 9443 12665 9495
rect 12717 9443 12755 9495
rect 12627 9402 12755 9443
rect 11494 9264 11622 9305
rect 11494 9212 11532 9264
rect 11584 9212 11622 9264
rect 11494 9171 11622 9212
rect 11494 8788 11622 8829
rect 11494 8736 11532 8788
rect 11584 8736 11622 8788
rect 11494 8695 11622 8736
rect 12627 8557 12755 8598
rect 12627 8505 12665 8557
rect 12717 8505 12755 8557
rect 12627 8464 12755 8505
rect 17423 8448 17551 8489
rect 17423 8396 17461 8448
rect 17513 8396 17551 8448
rect 17423 8355 17551 8396
rect 17800 7804 17928 7845
rect 17800 7752 17838 7804
rect 17890 7752 17928 7804
rect 12627 7695 12755 7736
rect 17800 7711 17928 7752
rect 12627 7643 12665 7695
rect 12717 7643 12755 7695
rect 12627 7602 12755 7643
rect 11494 7464 11622 7505
rect 11494 7412 11532 7464
rect 11584 7412 11622 7464
rect 11494 7371 11622 7412
rect 11494 6988 11622 7029
rect 11494 6936 11532 6988
rect 11584 6936 11622 6988
rect 11494 6895 11622 6936
rect 13004 6757 13132 6798
rect 13004 6705 13042 6757
rect 13094 6705 13132 6757
rect 13004 6664 13132 6705
rect 15156 6648 15284 6689
rect 15156 6596 15194 6648
rect 15246 6596 15284 6648
rect 15156 6555 15284 6596
rect 15534 6004 15662 6045
rect 15534 5952 15572 6004
rect 15624 5952 15662 6004
rect 13004 5895 13132 5936
rect 15534 5911 15662 5952
rect 13004 5843 13042 5895
rect 13094 5843 13132 5895
rect 13004 5802 13132 5843
rect 11494 5664 11622 5705
rect 11494 5612 11532 5664
rect 11584 5612 11622 5664
rect 11494 5571 11622 5612
rect 11494 5188 11622 5229
rect 11494 5136 11532 5188
rect 11584 5136 11622 5188
rect 11494 5095 11622 5136
rect 13004 4957 13132 4998
rect 13004 4905 13042 4957
rect 13094 4905 13132 4957
rect 13004 4864 13132 4905
rect 15912 4848 16040 4889
rect 15912 4796 15950 4848
rect 16002 4796 16040 4848
rect 15912 4755 16040 4796
rect 16290 4204 16418 4245
rect 16290 4152 16328 4204
rect 16380 4152 16418 4204
rect 13004 4095 13132 4136
rect 16290 4111 16418 4152
rect 13004 4043 13042 4095
rect 13094 4043 13132 4095
rect 13004 4002 13132 4043
rect 11494 3864 11622 3905
rect 11494 3812 11532 3864
rect 11584 3812 11622 3864
rect 11494 3771 11622 3812
rect 11494 3388 11622 3429
rect 11494 3336 11532 3388
rect 11584 3336 11622 3388
rect 11494 3295 11622 3336
rect 13004 3157 13132 3198
rect 13004 3105 13042 3157
rect 13094 3105 13132 3157
rect 13004 3064 13132 3105
rect 16667 3048 16795 3089
rect 16667 2996 16705 3048
rect 16757 2996 16795 3048
rect 16667 2955 16795 2996
rect 17045 2404 17173 2445
rect 17045 2352 17083 2404
rect 17135 2352 17173 2404
rect 13004 2295 13132 2336
rect 17045 2311 17173 2352
rect 13004 2243 13042 2295
rect 13094 2243 13132 2295
rect 13004 2202 13132 2243
rect 11494 2064 11622 2105
rect 11494 2012 11532 2064
rect 11584 2012 11622 2064
rect 11494 1971 11622 2012
rect 11494 1588 11622 1629
rect 11494 1536 11532 1588
rect 11584 1536 11622 1588
rect 11494 1495 11622 1536
rect 13004 1357 13132 1398
rect 13004 1305 13042 1357
rect 13094 1305 13132 1357
rect 13004 1264 13132 1305
rect 17423 1248 17551 1289
rect 17423 1196 17461 1248
rect 17513 1196 17551 1248
rect 17423 1155 17551 1196
rect 17800 604 17928 645
rect 17800 552 17838 604
rect 17890 552 17928 604
rect 13004 495 13132 536
rect 17800 511 17928 552
rect 13004 443 13042 495
rect 13094 443 13132 495
rect 13004 402 13132 443
rect 11493 264 11622 305
rect 11493 212 11532 264
rect 11584 212 11622 264
rect 11493 171 11622 212
rect 11871 171 12000 305
rect 12248 171 12378 305
rect 12626 171 12755 305
rect 13004 171 13133 305
rect 15156 171 15285 305
rect 15534 171 15663 305
rect 15911 171 16041 305
rect 16289 171 16418 305
rect 16667 171 16796 305
rect 17044 171 17174 305
rect 17422 171 17551 305
rect 17800 171 17929 305
rect 6835 -21 6965 112
<< metal3 >>
rect 765 13893 895 14027
rect 23358 13893 23487 14027
rect 765 12973 895 13107
rect 23358 12973 23487 13107
rect 765 12093 895 12227
rect 23358 12093 23487 12227
rect 765 11173 895 11307
rect 23358 11173 23487 11307
rect 765 10293 895 10427
rect 23358 10293 23487 10427
rect 765 9373 895 9507
rect 23358 9373 23487 9507
rect 765 8493 895 8627
rect 23358 8493 23487 8627
rect 765 7573 895 7707
rect 23358 7573 23487 7707
rect 765 6693 895 6827
rect 23358 6693 23487 6827
rect 765 5773 895 5907
rect 23358 5773 23487 5907
rect 765 4893 895 5027
rect 23358 4893 23487 5027
rect 765 3973 895 4107
rect 23358 3973 23487 4107
rect 765 3093 895 3227
rect 23358 3093 23487 3227
rect 765 2173 895 2307
rect 23358 2173 23487 2307
rect 765 1293 895 1427
rect 23358 1293 23487 1427
rect 765 373 895 507
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_0
timestamp 1666464484
transform 1 0 11558 0 1 1562
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_1
timestamp 1666464484
transform 1 0 11558 0 1 2038
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_2
timestamp 1666464484
transform 1 0 12691 0 1 7669
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_3
timestamp 1666464484
transform 1 0 12691 0 1 8531
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_4
timestamp 1666464484
transform 1 0 12691 0 1 9469
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_5
timestamp 1666464484
transform 1 0 12691 0 1 10331
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_6
timestamp 1666464484
transform 1 0 12691 0 1 11269
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_7
timestamp 1666464484
transform 1 0 12691 0 1 12131
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_8
timestamp 1666464484
transform 1 0 11558 0 1 14162
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_9
timestamp 1666464484
transform 1 0 11558 0 1 12362
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_10
timestamp 1666464484
transform 1 0 11558 0 1 10562
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_11
timestamp 1666464484
transform 1 0 11558 0 1 8762
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_12
timestamp 1666464484
transform 1 0 11558 0 1 6962
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_13
timestamp 1666464484
transform 1 0 11558 0 1 5162
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_14
timestamp 1666464484
transform 1 0 11558 0 1 3362
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_15
timestamp 1666464484
transform 1 0 13068 0 1 6731
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_16
timestamp 1666464484
transform 1 0 12691 0 1 13931
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_17
timestamp 1666464484
transform 1 0 12691 0 1 13069
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_18
timestamp 1666464484
transform 1 0 13068 0 1 469
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_19
timestamp 1666464484
transform 1 0 13068 0 1 1331
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_20
timestamp 1666464484
transform 1 0 13068 0 1 2269
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_21
timestamp 1666464484
transform 1 0 13068 0 1 3131
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_22
timestamp 1666464484
transform 1 0 13068 0 1 4069
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_23
timestamp 1666464484
transform 1 0 13068 0 1 4931
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_24
timestamp 1666464484
transform 1 0 13068 0 1 5869
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_25
timestamp 1666464484
transform 1 0 11558 0 1 12838
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_26
timestamp 1666464484
transform 1 0 11558 0 1 11038
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_27
timestamp 1666464484
transform 1 0 11558 0 1 9238
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_28
timestamp 1666464484
transform 1 0 11558 0 1 7438
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_29
timestamp 1666464484
transform 1 0 11558 0 1 5638
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_30
timestamp 1666464484
transform 1 0 11558 0 1 3838
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_31
timestamp 1666464484
transform 1 0 17864 0 1 578
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_32
timestamp 1666464484
transform 1 0 17487 0 1 1222
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_33
timestamp 1666464484
transform 1 0 17109 0 1 2378
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_34
timestamp 1666464484
transform 1 0 16731 0 1 3022
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_35
timestamp 1666464484
transform 1 0 16354 0 1 4178
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_36
timestamp 1666464484
transform 1 0 15976 0 1 4822
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_37
timestamp 1666464484
transform 1 0 15598 0 1 5978
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_38
timestamp 1666464484
transform 1 0 15220 0 1 6622
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_39
timestamp 1666464484
transform 1 0 15220 0 1 13822
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_40
timestamp 1666464484
transform 1 0 15598 0 1 13178
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_41
timestamp 1666464484
transform 1 0 15976 0 1 12022
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_42
timestamp 1666464484
transform 1 0 16354 0 1 11378
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_43
timestamp 1666464484
transform 1 0 16731 0 1 10222
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_44
timestamp 1666464484
transform 1 0 17109 0 1 9578
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_45
timestamp 1666464484
transform 1 0 17487 0 1 8422
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_46
timestamp 1666464484
transform 1 0 17864 0 1 7778
box 0 0 1 1
use M2_M1$$202394668_128x8m81  M2_M1$$202394668_128x8m81_47
timestamp 1666464484
transform 1 0 11558 0 1 238
box 0 0 1 1
use xdec8_128x8m81  xdec8_128x8m81_0
timestamp 1666464484
transform 1 0 0 0 1 7200
box 0 -228 24219 7428
use xdec8_128x8m81  xdec8_128x8m81_1
timestamp 1666464484
transform 1 0 0 0 1 0
box 0 -228 24219 7428
<< labels >>
rlabel metal3 s 830 5840 830 5840 4 LWL[6]
port 1 nsew
rlabel metal3 s 830 6760 830 6760 4 LWL[7]
port 2 nsew
rlabel metal3 s 23423 13960 23423 13960 4 RWL[15]
port 3 nsew
rlabel metal3 s 23423 13040 23423 13040 4 RWL[14]
port 4 nsew
rlabel metal3 s 23423 12160 23423 12160 4 RWL[13]
port 5 nsew
rlabel metal3 s 23423 11240 23423 11240 4 RWL[12]
port 6 nsew
rlabel metal3 s 830 8560 830 8560 4 LWL[9]
port 7 nsew
rlabel metal3 s 830 7640 830 7640 4 LWL[8]
port 8 nsew
rlabel metal3 s 830 440 830 440 4 LWL[0]
port 9 nsew
rlabel metal3 s 830 1360 830 1360 4 LWL[1]
port 10 nsew
rlabel metal3 s 830 2240 830 2240 4 LWL[2]
port 11 nsew
rlabel metal3 s 830 3160 830 3160 4 LWL[3]
port 12 nsew
rlabel metal3 s 830 4040 830 4040 4 LWL[4]
port 13 nsew
rlabel metal3 s 830 4960 830 4960 4 LWL[5]
port 14 nsew
rlabel metal3 s 23423 10360 23423 10360 4 RWL[11]
port 15 nsew
rlabel metal3 s 23423 9440 23423 9440 4 RWL[10]
port 16 nsew
rlabel metal3 s 23423 8560 23423 8560 4 RWL[9]
port 17 nsew
rlabel metal3 s 23423 7640 23423 7640 4 RWL[8]
port 18 nsew
rlabel metal3 s 23423 6760 23423 6760 4 RWL[7]
port 19 nsew
rlabel metal3 s 23423 4960 23423 4960 4 RWL[5]
port 20 nsew
rlabel metal3 s 23423 3160 23423 3160 4 RWL[3]
port 21 nsew
rlabel metal3 s 23423 1360 23423 1360 4 RWL[1]
port 22 nsew
rlabel metal3 s 23423 440 23423 440 4 RWL[0]
port 23 nsew
rlabel metal3 s 23423 2240 23423 2240 4 RWL[2]
port 24 nsew
rlabel metal3 s 830 13960 830 13960 4 LWL[15]
port 25 nsew
rlabel metal3 s 830 13040 830 13040 4 LWL[14]
port 26 nsew
rlabel metal3 s 830 12160 830 12160 4 LWL[13]
port 27 nsew
rlabel metal3 s 830 11240 830 11240 4 LWL[12]
port 28 nsew
rlabel metal3 s 830 10360 830 10360 4 LWL[11]
port 29 nsew
rlabel metal3 s 830 9440 830 9440 4 LWL[10]
port 30 nsew
rlabel metal3 s 23423 4040 23423 4040 4 RWL[4]
port 31 nsew
rlabel metal3 s 23423 5840 23423 5840 4 RWL[6]
port 32 nsew
rlabel metal2 s 17109 238 17109 238 4 xa[2]
port 33 nsew
rlabel metal2 s 6900 45 6900 45 4 men
port 34 nsew
rlabel metal2 s 17864 238 17864 238 4 xa[0]
port 35 nsew
rlabel metal2 s 16731 238 16731 238 4 xa[3]
port 36 nsew
rlabel metal2 s 16354 238 16354 238 4 xa[4]
port 37 nsew
rlabel metal2 s 15976 238 15976 238 4 xa[5]
port 38 nsew
rlabel metal2 s 15598 238 15598 238 4 xa[6]
port 39 nsew
rlabel metal2 s 15220 238 15220 238 4 xa[7]
port 40 nsew
rlabel metal2 s 11935 238 11935 238 4 xb[3]
port 41 nsew
rlabel metal2 s 12313 238 12313 238 4 xb[2]
port 42 nsew
rlabel metal2 s 12691 238 12691 238 4 xb[1]
port 43 nsew
rlabel metal2 s 13068 238 13068 238 4 xb[0]
port 44 nsew
rlabel metal2 s 11558 238 11558 238 4 xc
port 45 nsew
rlabel metal2 s 17487 238 17487 238 4 xa[1]
port 46 nsew
<< properties >>
string GDS_END 1698846
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1691536
<< end >>
