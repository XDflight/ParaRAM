magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 148 75 312 1728
<< metal2 >>
rect 360 0 460 1405
<< metal3 >>
rect -511 630 489 2425
rect 714 1817 1714 2425
use M2_M14310590548783_128x8m81  M2_M14310590548783_128x8m81_0
timestamp 1666464484
transform 1 0 1214 0 1 1981
box -472 -162 472 162
use M3_M24310590548776_128x8m81  M3_M24310590548776_128x8m81_0
timestamp 1666464484
transform 1 0 1214 0 1 1981
box -472 -162 472 162
use M3_M24310590548781_128x8m81  M3_M24310590548781_128x8m81_0
timestamp 1666464484
transform 1 0 -12 0 1 1126
box -472 -472 472 472
<< properties >>
string GDS_END 1485964
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 1485578
string path -0.055 3.150 -0.055 12.125 
<< end >>
