magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect 0 69946 1000 69968
rect 0 69897 177 69946
rect 0 13151 25 69897
rect 71 69800 177 69897
rect 823 69897 1000 69946
rect 823 69800 929 69897
rect 71 69778 929 69800
rect 71 13287 93 69778
rect 907 13287 929 69778
rect 71 13265 929 13287
rect 71 13151 177 13265
rect 0 13119 177 13151
rect 823 13151 929 13265
rect 975 13151 1000 69897
rect 823 13119 1000 13151
rect 0 13097 1000 13119
<< psubdiffcont >>
rect 25 13151 71 69897
rect 177 69800 823 69946
rect 177 13119 823 13265
rect 929 13151 975 69897
<< metal1 >>
rect -32 69946 1032 69957
rect -32 69897 177 69946
rect -32 13151 25 69897
rect 71 69800 177 69897
rect 823 69897 1032 69946
rect 823 69800 929 69897
rect 71 69789 929 69800
rect 71 64896 82 69789
rect 71 64884 123 64896
rect 111 64832 123 64884
rect 71 64760 123 64832
rect 111 64708 123 64760
rect 71 64636 123 64708
rect 111 64584 123 64636
rect 71 64512 123 64584
rect 111 64460 123 64512
rect 71 64388 123 64460
rect 111 64336 123 64388
rect 71 64264 123 64336
rect 111 64212 123 64264
rect 71 64140 123 64212
rect 111 64088 123 64140
rect 71 64016 123 64088
rect 111 63964 123 64016
rect 71 63892 123 63964
rect 111 63840 123 63892
rect 71 63768 123 63840
rect 111 63716 123 63768
rect 71 63704 123 63716
rect 839 64884 915 64896
rect 839 64832 851 64884
rect 903 64832 915 64884
rect 839 64760 915 64832
rect 839 64708 851 64760
rect 903 64708 915 64760
rect 839 64636 915 64708
rect 839 64584 851 64636
rect 903 64584 915 64636
rect 839 64512 915 64584
rect 839 64460 851 64512
rect 903 64460 915 64512
rect 839 64388 915 64460
rect 839 64336 851 64388
rect 903 64336 915 64388
rect 839 64264 915 64336
rect 839 64212 851 64264
rect 903 64212 915 64264
rect 839 64140 915 64212
rect 839 64088 851 64140
rect 903 64088 915 64140
rect 839 64016 915 64088
rect 839 63964 851 64016
rect 903 63964 915 64016
rect 839 63892 915 63964
rect 839 63840 851 63892
rect 903 63840 915 63892
rect 839 63768 915 63840
rect 839 63716 851 63768
rect 903 63716 915 63768
rect 839 63704 915 63716
rect 71 50496 82 63704
rect 71 50484 123 50496
rect 111 50432 123 50484
rect 71 50360 123 50432
rect 111 50308 123 50360
rect 71 50236 123 50308
rect 111 50184 123 50236
rect 71 50112 123 50184
rect 111 50060 123 50112
rect 71 49988 123 50060
rect 111 49936 123 49988
rect 71 49864 123 49936
rect 111 49812 123 49864
rect 71 49740 123 49812
rect 111 49688 123 49740
rect 71 49616 123 49688
rect 111 49564 123 49616
rect 71 49492 123 49564
rect 111 49440 123 49492
rect 71 49368 123 49440
rect 111 49316 123 49368
rect 71 49304 123 49316
rect 839 50484 915 50496
rect 839 50432 851 50484
rect 903 50432 915 50484
rect 839 50360 915 50432
rect 839 50308 851 50360
rect 903 50308 915 50360
rect 839 50236 915 50308
rect 839 50184 851 50236
rect 903 50184 915 50236
rect 839 50112 915 50184
rect 839 50060 851 50112
rect 903 50060 915 50112
rect 839 49988 915 50060
rect 839 49936 851 49988
rect 903 49936 915 49988
rect 839 49864 915 49936
rect 839 49812 851 49864
rect 903 49812 915 49864
rect 839 49740 915 49812
rect 839 49688 851 49740
rect 903 49688 915 49740
rect 839 49616 915 49688
rect 839 49564 851 49616
rect 903 49564 915 49616
rect 839 49492 915 49564
rect 839 49440 851 49492
rect 903 49440 915 49492
rect 839 49368 915 49440
rect 839 49316 851 49368
rect 903 49316 915 49368
rect 839 49304 915 49316
rect 71 13276 82 49304
rect 918 13276 929 69789
rect 71 13265 929 13276
rect 71 13151 177 13265
rect -32 13119 177 13151
rect 823 13151 929 13265
rect 975 13151 1032 69897
rect 823 13119 1032 13151
rect -32 13108 1032 13119
<< via1 >>
rect 59 64832 71 64884
rect 71 64832 111 64884
rect 59 64708 71 64760
rect 71 64708 111 64760
rect 59 64584 71 64636
rect 71 64584 111 64636
rect 59 64460 71 64512
rect 71 64460 111 64512
rect 59 64336 71 64388
rect 71 64336 111 64388
rect 59 64212 71 64264
rect 71 64212 111 64264
rect 59 64088 71 64140
rect 71 64088 111 64140
rect 59 63964 71 64016
rect 71 63964 111 64016
rect 59 63840 71 63892
rect 71 63840 111 63892
rect 59 63716 71 63768
rect 71 63716 111 63768
rect 851 64832 903 64884
rect 851 64708 903 64760
rect 851 64584 903 64636
rect 851 64460 903 64512
rect 851 64336 903 64388
rect 851 64212 903 64264
rect 851 64088 903 64140
rect 851 63964 903 64016
rect 851 63840 903 63892
rect 851 63716 903 63768
rect 59 50432 71 50484
rect 71 50432 111 50484
rect 59 50308 71 50360
rect 71 50308 111 50360
rect 59 50184 71 50236
rect 71 50184 111 50236
rect 59 50060 71 50112
rect 71 50060 111 50112
rect 59 49936 71 49988
rect 71 49936 111 49988
rect 59 49812 71 49864
rect 71 49812 111 49864
rect 59 49688 71 49740
rect 71 49688 111 49740
rect 59 49564 71 49616
rect 71 49564 111 49616
rect 59 49440 71 49492
rect 71 49440 111 49492
rect 59 49316 71 49368
rect 71 49316 111 49368
rect 851 50432 903 50484
rect 851 50308 903 50360
rect 851 50184 903 50236
rect 851 50060 903 50112
rect 851 49936 903 49988
rect 851 49812 903 49864
rect 851 49688 903 49740
rect 851 49564 903 49616
rect 851 49440 903 49492
rect 851 49316 903 49368
<< metal2 >>
rect 56 65000 178 69660
rect 656 69579 732 69589
rect 656 69523 666 69579
rect 722 69523 732 69579
rect 656 69447 732 69523
rect 656 69391 666 69447
rect 722 69391 732 69447
rect 656 69315 732 69391
rect 656 69259 666 69315
rect 722 69259 732 69315
rect 656 69183 732 69259
rect 656 69127 666 69183
rect 722 69127 732 69183
rect 656 69051 732 69127
rect 656 68995 666 69051
rect 722 68995 732 69051
rect 656 68919 732 68995
rect 656 68863 666 68919
rect 722 68863 732 68919
rect 656 68787 732 68863
rect 656 68731 666 68787
rect 722 68731 732 68787
rect 656 68655 732 68731
rect 656 68599 666 68655
rect 722 68599 732 68655
rect 656 68523 732 68599
rect 656 68467 666 68523
rect 722 68467 732 68523
rect 0 64886 178 65000
rect 0 64830 57 64886
rect 113 64830 178 64886
rect 0 64762 178 64830
rect 0 64706 57 64762
rect 113 64706 178 64762
rect 0 64638 178 64706
rect 0 64582 57 64638
rect 113 64582 178 64638
rect 0 64514 178 64582
rect 0 64458 57 64514
rect 113 64458 178 64514
rect 0 64390 178 64458
rect 0 64334 57 64390
rect 113 64334 178 64390
rect 0 64266 178 64334
rect 0 64210 57 64266
rect 113 64210 178 64266
rect 0 64142 178 64210
rect 0 64086 57 64142
rect 113 64086 178 64142
rect 0 64018 178 64086
rect 0 63962 57 64018
rect 113 63962 178 64018
rect 0 63894 178 63962
rect 0 63838 57 63894
rect 113 63838 178 63894
rect 0 63770 178 63838
rect 0 63714 57 63770
rect 113 63714 178 63770
rect 0 63600 178 63714
rect 56 50600 178 63600
rect 0 50486 178 50600
rect 0 50430 57 50486
rect 113 50430 178 50486
rect 0 50362 178 50430
rect 0 50306 57 50362
rect 113 50306 178 50362
rect 0 50238 178 50306
rect 0 50182 57 50238
rect 113 50182 178 50238
rect 0 50114 178 50182
rect 0 50058 57 50114
rect 113 50058 178 50114
rect 0 49990 178 50058
rect 0 49934 57 49990
rect 113 49934 178 49990
rect 0 49866 178 49934
rect 0 49810 57 49866
rect 113 49810 178 49866
rect 0 49742 178 49810
rect 0 49686 57 49742
rect 113 49686 178 49742
rect 0 49618 178 49686
rect 0 49562 57 49618
rect 113 49562 178 49618
rect 0 49494 178 49562
rect 0 49438 57 49494
rect 113 49438 178 49494
rect 0 49370 178 49438
rect 0 49314 57 49370
rect 113 49314 178 49370
rect 0 49200 178 49314
rect 56 13491 178 49200
rect 280 68050 356 68189
rect 280 67994 290 68050
rect 346 67994 356 68050
rect 280 67918 356 67994
rect 280 67862 290 67918
rect 346 67862 356 67918
rect 280 67786 356 67862
rect 280 67730 290 67786
rect 346 67730 356 67786
rect 280 67654 356 67730
rect 280 67598 290 67654
rect 346 67598 356 67654
rect 280 67522 356 67598
rect 280 67466 290 67522
rect 346 67466 356 67522
rect 280 67390 356 67466
rect 280 67334 290 67390
rect 346 67334 356 67390
rect 280 67258 356 67334
rect 280 67202 290 67258
rect 346 67202 356 67258
rect 280 67126 356 67202
rect 280 67070 290 67126
rect 346 67070 356 67126
rect 280 66994 356 67070
rect 280 66938 290 66994
rect 346 66938 356 66994
rect 280 60061 356 66938
rect 656 66466 732 68467
rect 656 66410 666 66466
rect 722 66410 732 66466
rect 656 66334 732 66410
rect 656 66278 666 66334
rect 722 66278 732 66334
rect 656 66202 732 66278
rect 656 66146 666 66202
rect 722 66146 732 66202
rect 656 66070 732 66146
rect 656 66014 666 66070
rect 722 66014 732 66070
rect 656 65938 732 66014
rect 656 65882 666 65938
rect 722 65882 732 65938
rect 656 65806 732 65882
rect 656 65750 666 65806
rect 722 65750 732 65806
rect 656 65674 732 65750
rect 656 65618 666 65674
rect 722 65618 732 65674
rect 656 65542 732 65618
rect 656 65486 666 65542
rect 722 65486 732 65542
rect 656 65410 732 65486
rect 656 65354 666 65410
rect 722 65354 732 65410
rect 472 63253 548 63263
rect 472 63197 482 63253
rect 538 63197 548 63253
rect 472 63121 548 63197
rect 472 63065 482 63121
rect 538 63065 548 63121
rect 472 62989 548 63065
rect 472 62933 482 62989
rect 538 62933 548 62989
rect 472 62857 548 62933
rect 472 62801 482 62857
rect 538 62801 548 62857
rect 472 62725 548 62801
rect 472 62669 482 62725
rect 538 62669 548 62725
rect 472 62593 548 62669
rect 472 62537 482 62593
rect 538 62537 548 62593
rect 472 62461 548 62537
rect 472 62405 482 62461
rect 538 62405 548 62461
rect 472 62329 548 62405
rect 472 62273 482 62329
rect 538 62273 548 62329
rect 472 62197 548 62273
rect 472 62141 482 62197
rect 538 62141 548 62197
rect 472 62131 548 62141
rect 280 60005 290 60061
rect 346 60005 356 60061
rect 280 59929 356 60005
rect 280 59873 290 59929
rect 346 59873 356 59929
rect 280 59797 356 59873
rect 280 59741 290 59797
rect 346 59741 356 59797
rect 280 59665 356 59741
rect 280 59609 290 59665
rect 346 59609 356 59665
rect 280 59533 356 59609
rect 280 59477 290 59533
rect 346 59477 356 59533
rect 280 59401 356 59477
rect 280 59345 290 59401
rect 346 59345 356 59401
rect 280 59269 356 59345
rect 280 59213 290 59269
rect 346 59213 356 59269
rect 280 59137 356 59213
rect 280 59081 290 59137
rect 346 59081 356 59137
rect 280 59005 356 59081
rect 280 58949 290 59005
rect 346 58949 356 59005
rect 280 56879 356 58949
rect 280 56823 290 56879
rect 346 56823 356 56879
rect 280 56747 356 56823
rect 280 56691 290 56747
rect 346 56691 356 56747
rect 280 56615 356 56691
rect 280 56559 290 56615
rect 346 56559 356 56615
rect 280 56483 356 56559
rect 280 56427 290 56483
rect 346 56427 356 56483
rect 280 56351 356 56427
rect 280 56295 290 56351
rect 346 56295 356 56351
rect 280 56219 356 56295
rect 280 56163 290 56219
rect 346 56163 356 56219
rect 280 56087 356 56163
rect 280 56031 290 56087
rect 346 56031 356 56087
rect 280 55955 356 56031
rect 280 55899 290 55955
rect 346 55899 356 55955
rect 280 55823 356 55899
rect 280 55767 290 55823
rect 346 55767 356 55823
rect 280 55260 356 55767
rect 280 55204 290 55260
rect 346 55204 356 55260
rect 280 55128 356 55204
rect 280 55072 290 55128
rect 346 55072 356 55128
rect 280 54996 356 55072
rect 280 54940 290 54996
rect 346 54940 356 54996
rect 280 54864 356 54940
rect 280 54808 290 54864
rect 346 54808 356 54864
rect 280 54732 356 54808
rect 280 54676 290 54732
rect 346 54676 356 54732
rect 280 54600 356 54676
rect 280 54544 290 54600
rect 346 54544 356 54600
rect 280 54468 356 54544
rect 280 54412 290 54468
rect 346 54412 356 54468
rect 280 54336 356 54412
rect 280 54280 290 54336
rect 346 54280 356 54336
rect 280 54204 356 54280
rect 280 54148 290 54204
rect 346 54148 356 54204
rect 280 53669 356 54148
rect 280 53613 290 53669
rect 346 53613 356 53669
rect 280 53537 356 53613
rect 280 53481 290 53537
rect 346 53481 356 53537
rect 280 53405 356 53481
rect 280 53349 290 53405
rect 346 53349 356 53405
rect 280 53273 356 53349
rect 280 53217 290 53273
rect 346 53217 356 53273
rect 280 53141 356 53217
rect 280 53085 290 53141
rect 346 53085 356 53141
rect 280 53009 356 53085
rect 280 52953 290 53009
rect 346 52953 356 53009
rect 280 52877 356 52953
rect 280 52821 290 52877
rect 346 52821 356 52877
rect 280 52745 356 52821
rect 280 52689 290 52745
rect 346 52689 356 52745
rect 280 52613 356 52689
rect 280 52557 290 52613
rect 346 52557 356 52613
rect 280 45593 356 52557
rect 656 61664 732 65354
rect 656 61608 666 61664
rect 722 61608 732 61664
rect 656 61532 732 61608
rect 656 61476 666 61532
rect 722 61476 732 61532
rect 656 61400 732 61476
rect 656 61344 666 61400
rect 722 61344 732 61400
rect 656 61268 732 61344
rect 656 61212 666 61268
rect 722 61212 732 61268
rect 656 61136 732 61212
rect 656 61080 666 61136
rect 722 61080 732 61136
rect 656 61004 732 61080
rect 656 60948 666 61004
rect 722 60948 732 61004
rect 656 60872 732 60948
rect 656 60816 666 60872
rect 722 60816 732 60872
rect 656 60740 732 60816
rect 656 60684 666 60740
rect 722 60684 732 60740
rect 656 60608 732 60684
rect 656 60552 666 60608
rect 722 60552 732 60608
rect 656 58453 732 60552
rect 656 58397 666 58453
rect 722 58397 732 58453
rect 656 58321 732 58397
rect 656 58265 666 58321
rect 722 58265 732 58321
rect 656 58189 732 58265
rect 656 58133 666 58189
rect 722 58133 732 58189
rect 656 58057 732 58133
rect 656 58001 666 58057
rect 722 58001 732 58057
rect 656 57925 732 58001
rect 656 57869 666 57925
rect 722 57869 732 57925
rect 656 57793 732 57869
rect 656 57737 666 57793
rect 722 57737 732 57793
rect 656 57661 732 57737
rect 656 57605 666 57661
rect 722 57605 732 57661
rect 656 57529 732 57605
rect 656 57473 666 57529
rect 722 57473 732 57529
rect 656 57397 732 57473
rect 656 57341 666 57397
rect 722 57341 732 57397
rect 472 52060 548 52070
rect 472 52004 482 52060
rect 538 52004 548 52060
rect 472 51928 548 52004
rect 472 51872 482 51928
rect 538 51872 548 51928
rect 472 51796 548 51872
rect 472 51740 482 51796
rect 538 51740 548 51796
rect 472 51664 548 51740
rect 472 51608 482 51664
rect 538 51608 548 51664
rect 472 51532 548 51608
rect 472 51476 482 51532
rect 538 51476 548 51532
rect 472 51400 548 51476
rect 472 51344 482 51400
rect 538 51344 548 51400
rect 472 51268 548 51344
rect 472 51212 482 51268
rect 538 51212 548 51268
rect 472 51136 548 51212
rect 472 51080 482 51136
rect 538 51080 548 51136
rect 472 51004 548 51080
rect 472 50948 482 51004
rect 538 50948 548 51004
rect 472 50938 548 50948
rect 280 45537 290 45593
rect 346 45537 356 45593
rect 280 45461 356 45537
rect 280 45405 290 45461
rect 346 45405 356 45461
rect 280 45329 356 45405
rect 280 45273 290 45329
rect 346 45273 356 45329
rect 280 45197 356 45273
rect 280 45141 290 45197
rect 346 45141 356 45197
rect 280 45065 356 45141
rect 280 45009 290 45065
rect 346 45009 356 45065
rect 280 44933 356 45009
rect 280 44877 290 44933
rect 346 44877 356 44933
rect 280 44801 356 44877
rect 280 44745 290 44801
rect 346 44745 356 44801
rect 280 44669 356 44745
rect 280 44613 290 44669
rect 346 44613 356 44669
rect 280 44537 356 44613
rect 280 44481 290 44537
rect 346 44481 356 44537
rect 280 44405 356 44481
rect 280 44349 290 44405
rect 346 44349 356 44405
rect 280 44273 356 44349
rect 280 44217 290 44273
rect 346 44217 356 44273
rect 280 44141 356 44217
rect 280 44085 290 44141
rect 346 44085 356 44141
rect 280 44009 356 44085
rect 280 43953 290 44009
rect 346 43953 356 44009
rect 280 43877 356 43953
rect 280 43821 290 43877
rect 346 43821 356 43877
rect 280 43745 356 43821
rect 280 43689 290 43745
rect 346 43689 356 43745
rect 280 43613 356 43689
rect 280 43557 290 43613
rect 346 43557 356 43613
rect 280 43481 356 43557
rect 280 43425 290 43481
rect 346 43425 356 43481
rect 280 43349 356 43425
rect 280 43293 290 43349
rect 346 43293 356 43349
rect 280 43217 356 43293
rect 280 43161 290 43217
rect 346 43161 356 43217
rect 280 43085 356 43161
rect 280 43029 290 43085
rect 346 43029 356 43085
rect 280 42451 356 43029
rect 280 42395 290 42451
rect 346 42395 356 42451
rect 280 42319 356 42395
rect 280 42263 290 42319
rect 346 42263 356 42319
rect 280 42187 356 42263
rect 280 42131 290 42187
rect 346 42131 356 42187
rect 280 42055 356 42131
rect 280 41999 290 42055
rect 346 41999 356 42055
rect 280 41923 356 41999
rect 280 41867 290 41923
rect 346 41867 356 41923
rect 280 41791 356 41867
rect 280 41735 290 41791
rect 346 41735 356 41791
rect 280 41659 356 41735
rect 280 41603 290 41659
rect 346 41603 356 41659
rect 280 41527 356 41603
rect 280 41471 290 41527
rect 346 41471 356 41527
rect 280 41395 356 41471
rect 280 41339 290 41395
rect 346 41339 356 41395
rect 280 39170 356 41339
rect 280 39114 290 39170
rect 346 39114 356 39170
rect 280 39038 356 39114
rect 280 38982 290 39038
rect 346 38982 356 39038
rect 280 38906 356 38982
rect 280 38850 290 38906
rect 346 38850 356 38906
rect 280 38774 356 38850
rect 280 38718 290 38774
rect 346 38718 356 38774
rect 280 38642 356 38718
rect 280 38586 290 38642
rect 346 38586 356 38642
rect 280 38510 356 38586
rect 280 38454 290 38510
rect 346 38454 356 38510
rect 280 38378 356 38454
rect 280 38322 290 38378
rect 346 38322 356 38378
rect 280 38246 356 38322
rect 280 38190 290 38246
rect 346 38190 356 38246
rect 280 38114 356 38190
rect 280 38058 290 38114
rect 346 38058 356 38114
rect 280 37982 356 38058
rect 280 37926 290 37982
rect 346 37926 356 37982
rect 280 37850 356 37926
rect 280 37794 290 37850
rect 346 37794 356 37850
rect 280 37718 356 37794
rect 280 37662 290 37718
rect 346 37662 356 37718
rect 280 37586 356 37662
rect 280 37530 290 37586
rect 346 37530 356 37586
rect 280 37454 356 37530
rect 280 37398 290 37454
rect 346 37398 356 37454
rect 280 37322 356 37398
rect 280 37266 290 37322
rect 346 37266 356 37322
rect 280 37190 356 37266
rect 280 37134 290 37190
rect 346 37134 356 37190
rect 280 37058 356 37134
rect 280 37002 290 37058
rect 346 37002 356 37058
rect 280 36926 356 37002
rect 280 36870 290 36926
rect 346 36870 356 36926
rect 280 36794 356 36870
rect 280 36738 290 36794
rect 346 36738 356 36794
rect 280 36662 356 36738
rect 280 36606 290 36662
rect 346 36606 356 36662
rect 280 36000 356 36606
rect 280 35944 290 36000
rect 346 35944 356 36000
rect 280 35868 356 35944
rect 280 35812 290 35868
rect 346 35812 356 35868
rect 280 35736 356 35812
rect 280 35680 290 35736
rect 346 35680 356 35736
rect 280 35604 356 35680
rect 280 35548 290 35604
rect 346 35548 356 35604
rect 280 35472 356 35548
rect 280 35416 290 35472
rect 346 35416 356 35472
rect 280 35340 356 35416
rect 280 35284 290 35340
rect 346 35284 356 35340
rect 280 35208 356 35284
rect 280 35152 290 35208
rect 346 35152 356 35208
rect 280 35076 356 35152
rect 280 35020 290 35076
rect 346 35020 356 35076
rect 280 34944 356 35020
rect 280 34888 290 34944
rect 346 34888 356 34944
rect 280 34812 356 34888
rect 280 34756 290 34812
rect 346 34756 356 34812
rect 280 34680 356 34756
rect 280 34624 290 34680
rect 346 34624 356 34680
rect 280 34548 356 34624
rect 280 34492 290 34548
rect 346 34492 356 34548
rect 280 34416 356 34492
rect 280 34360 290 34416
rect 346 34360 356 34416
rect 280 34284 356 34360
rect 280 34228 290 34284
rect 346 34228 356 34284
rect 280 34152 356 34228
rect 280 34096 290 34152
rect 346 34096 356 34152
rect 280 34020 356 34096
rect 280 33964 290 34020
rect 346 33964 356 34020
rect 280 33888 356 33964
rect 280 33832 290 33888
rect 346 33832 356 33888
rect 280 33756 356 33832
rect 280 33700 290 33756
rect 346 33700 356 33756
rect 280 33624 356 33700
rect 280 33568 290 33624
rect 346 33568 356 33624
rect 280 33492 356 33568
rect 280 33436 290 33492
rect 346 33436 356 33492
rect 280 32795 356 33436
rect 280 32739 290 32795
rect 346 32739 356 32795
rect 280 32663 356 32739
rect 280 32607 290 32663
rect 346 32607 356 32663
rect 280 32531 356 32607
rect 280 32475 290 32531
rect 346 32475 356 32531
rect 280 32399 356 32475
rect 280 32343 290 32399
rect 346 32343 356 32399
rect 280 32267 356 32343
rect 280 32211 290 32267
rect 346 32211 356 32267
rect 280 32135 356 32211
rect 280 32079 290 32135
rect 346 32079 356 32135
rect 280 32003 356 32079
rect 280 31947 290 32003
rect 346 31947 356 32003
rect 280 31871 356 31947
rect 280 31815 290 31871
rect 346 31815 356 31871
rect 280 31739 356 31815
rect 280 31683 290 31739
rect 346 31683 356 31739
rect 280 31607 356 31683
rect 280 31551 290 31607
rect 346 31551 356 31607
rect 280 31475 356 31551
rect 280 31419 290 31475
rect 346 31419 356 31475
rect 280 31343 356 31419
rect 280 31287 290 31343
rect 346 31287 356 31343
rect 280 31211 356 31287
rect 280 31155 290 31211
rect 346 31155 356 31211
rect 280 31079 356 31155
rect 280 31023 290 31079
rect 346 31023 356 31079
rect 280 30947 356 31023
rect 280 30891 290 30947
rect 346 30891 356 30947
rect 280 30815 356 30891
rect 280 30759 290 30815
rect 346 30759 356 30815
rect 280 30683 356 30759
rect 280 30627 290 30683
rect 346 30627 356 30683
rect 280 30551 356 30627
rect 280 30495 290 30551
rect 346 30495 356 30551
rect 280 30419 356 30495
rect 280 30363 290 30419
rect 346 30363 356 30419
rect 280 30287 356 30363
rect 280 30231 290 30287
rect 346 30231 356 30287
rect 280 29625 356 30231
rect 280 29569 290 29625
rect 346 29569 356 29625
rect 280 29493 356 29569
rect 280 29437 290 29493
rect 346 29437 356 29493
rect 280 29361 356 29437
rect 280 29305 290 29361
rect 346 29305 356 29361
rect 280 29229 356 29305
rect 280 29173 290 29229
rect 346 29173 356 29229
rect 280 29097 356 29173
rect 280 29041 290 29097
rect 346 29041 356 29097
rect 280 28965 356 29041
rect 280 28909 290 28965
rect 346 28909 356 28965
rect 280 28833 356 28909
rect 280 28777 290 28833
rect 346 28777 356 28833
rect 280 28701 356 28777
rect 280 28645 290 28701
rect 346 28645 356 28701
rect 280 28569 356 28645
rect 280 28513 290 28569
rect 346 28513 356 28569
rect 280 28437 356 28513
rect 280 28381 290 28437
rect 346 28381 356 28437
rect 280 28305 356 28381
rect 280 28249 290 28305
rect 346 28249 356 28305
rect 280 28173 356 28249
rect 280 28117 290 28173
rect 346 28117 356 28173
rect 280 28041 356 28117
rect 280 27985 290 28041
rect 346 27985 356 28041
rect 280 27909 356 27985
rect 280 27853 290 27909
rect 346 27853 356 27909
rect 280 27777 356 27853
rect 280 27721 290 27777
rect 346 27721 356 27777
rect 280 27645 356 27721
rect 280 27589 290 27645
rect 346 27589 356 27645
rect 280 27513 356 27589
rect 280 27457 290 27513
rect 346 27457 356 27513
rect 280 27381 356 27457
rect 280 27325 290 27381
rect 346 27325 356 27381
rect 280 27249 356 27325
rect 280 27193 290 27249
rect 346 27193 356 27249
rect 280 27117 356 27193
rect 280 27061 290 27117
rect 346 27061 356 27117
rect 280 24854 356 27061
rect 280 24798 290 24854
rect 346 24798 356 24854
rect 280 24722 356 24798
rect 280 24666 290 24722
rect 346 24666 356 24722
rect 280 24590 356 24666
rect 280 24534 290 24590
rect 346 24534 356 24590
rect 280 24458 356 24534
rect 280 24402 290 24458
rect 346 24402 356 24458
rect 280 24326 356 24402
rect 280 24270 290 24326
rect 346 24270 356 24326
rect 280 24194 356 24270
rect 280 24138 290 24194
rect 346 24138 356 24194
rect 280 24062 356 24138
rect 280 24006 290 24062
rect 346 24006 356 24062
rect 280 23930 356 24006
rect 280 23874 290 23930
rect 346 23874 356 23930
rect 280 23798 356 23874
rect 280 23742 290 23798
rect 346 23742 356 23798
rect 280 23600 356 23742
rect 656 48810 732 57341
rect 656 48754 666 48810
rect 722 48754 732 48810
rect 656 48678 732 48754
rect 656 48622 666 48678
rect 722 48622 732 48678
rect 656 48546 732 48622
rect 656 48490 666 48546
rect 722 48490 732 48546
rect 656 48414 732 48490
rect 656 48358 666 48414
rect 722 48358 732 48414
rect 656 48282 732 48358
rect 656 48226 666 48282
rect 722 48226 732 48282
rect 656 48150 732 48226
rect 656 48094 666 48150
rect 722 48094 732 48150
rect 656 48018 732 48094
rect 656 47962 666 48018
rect 722 47962 732 48018
rect 656 47886 732 47962
rect 656 47830 666 47886
rect 722 47830 732 47886
rect 656 47754 732 47830
rect 656 47698 666 47754
rect 722 47698 732 47754
rect 656 47622 732 47698
rect 656 47566 666 47622
rect 722 47566 732 47622
rect 656 47490 732 47566
rect 656 47434 666 47490
rect 722 47434 732 47490
rect 656 47358 732 47434
rect 656 47302 666 47358
rect 722 47302 732 47358
rect 656 47226 732 47302
rect 656 47170 666 47226
rect 722 47170 732 47226
rect 656 47094 732 47170
rect 656 47038 666 47094
rect 722 47038 732 47094
rect 656 46962 732 47038
rect 656 46906 666 46962
rect 722 46906 732 46962
rect 656 46830 732 46906
rect 656 46774 666 46830
rect 722 46774 732 46830
rect 656 46698 732 46774
rect 656 46642 666 46698
rect 722 46642 732 46698
rect 656 46566 732 46642
rect 656 46510 666 46566
rect 722 46510 732 46566
rect 656 46434 732 46510
rect 656 46378 666 46434
rect 722 46378 732 46434
rect 656 46302 732 46378
rect 656 46246 666 46302
rect 722 46246 732 46302
rect 656 40883 732 46246
rect 656 40827 666 40883
rect 722 40827 732 40883
rect 656 40751 732 40827
rect 656 40695 666 40751
rect 722 40695 732 40751
rect 656 40619 732 40695
rect 656 40563 666 40619
rect 722 40563 732 40619
rect 656 40487 732 40563
rect 656 40431 666 40487
rect 722 40431 732 40487
rect 656 40355 732 40431
rect 656 40299 666 40355
rect 722 40299 732 40355
rect 656 40223 732 40299
rect 656 40167 666 40223
rect 722 40167 732 40223
rect 656 40091 732 40167
rect 656 40035 666 40091
rect 722 40035 732 40091
rect 656 39959 732 40035
rect 656 39903 666 39959
rect 722 39903 732 39959
rect 656 39827 732 39903
rect 656 39771 666 39827
rect 722 39771 732 39827
rect 656 26485 732 39771
rect 656 26429 666 26485
rect 722 26429 732 26485
rect 656 26353 732 26429
rect 656 26297 666 26353
rect 722 26297 732 26353
rect 656 26221 732 26297
rect 656 26165 666 26221
rect 722 26165 732 26221
rect 656 26089 732 26165
rect 656 26033 666 26089
rect 722 26033 732 26089
rect 656 25957 732 26033
rect 656 25901 666 25957
rect 722 25901 732 25957
rect 656 25825 732 25901
rect 656 25769 666 25825
rect 722 25769 732 25825
rect 656 25693 732 25769
rect 656 25637 666 25693
rect 722 25637 732 25693
rect 656 25561 732 25637
rect 656 25505 666 25561
rect 722 25505 732 25561
rect 656 25429 732 25505
rect 656 25373 666 25429
rect 722 25373 732 25429
rect 656 23190 732 25373
rect 656 23134 666 23190
rect 722 23134 732 23190
rect 656 23058 732 23134
rect 656 23002 666 23058
rect 722 23002 732 23058
rect 656 22926 732 23002
rect 656 22870 666 22926
rect 722 22870 732 22926
rect 656 22794 732 22870
rect 656 22738 666 22794
rect 722 22738 732 22794
rect 656 22662 732 22738
rect 656 22606 666 22662
rect 722 22606 732 22662
rect 656 22530 732 22606
rect 656 22474 666 22530
rect 722 22474 732 22530
rect 656 22398 732 22474
rect 656 22342 666 22398
rect 722 22342 732 22398
rect 656 22266 732 22342
rect 656 22210 666 22266
rect 722 22210 732 22266
rect 656 22134 732 22210
rect 656 22078 666 22134
rect 722 22078 732 22134
rect 656 22002 732 22078
rect 656 21946 666 22002
rect 722 21946 732 22002
rect 656 21870 732 21946
rect 656 21814 666 21870
rect 722 21814 732 21870
rect 656 21738 732 21814
rect 656 21682 666 21738
rect 722 21682 732 21738
rect 656 21606 732 21682
rect 656 21550 666 21606
rect 722 21550 732 21606
rect 656 21474 732 21550
rect 656 21418 666 21474
rect 722 21418 732 21474
rect 656 21342 732 21418
rect 656 21286 666 21342
rect 722 21286 732 21342
rect 656 21210 732 21286
rect 656 21154 666 21210
rect 722 21154 732 21210
rect 656 21078 732 21154
rect 656 21022 666 21078
rect 722 21022 732 21078
rect 656 20946 732 21022
rect 656 20890 666 20946
rect 722 20890 732 20946
rect 656 20814 732 20890
rect 656 20758 666 20814
rect 722 20758 732 20814
rect 656 20682 732 20758
rect 656 20626 666 20682
rect 722 20626 732 20682
rect 656 19978 732 20626
rect 656 19922 666 19978
rect 722 19922 732 19978
rect 656 19846 732 19922
rect 656 19790 666 19846
rect 722 19790 732 19846
rect 656 19714 732 19790
rect 656 19658 666 19714
rect 722 19658 732 19714
rect 656 19582 732 19658
rect 656 19526 666 19582
rect 722 19526 732 19582
rect 656 19450 732 19526
rect 656 19394 666 19450
rect 722 19394 732 19450
rect 656 19318 732 19394
rect 656 19262 666 19318
rect 722 19262 732 19318
rect 656 19186 732 19262
rect 656 19130 666 19186
rect 722 19130 732 19186
rect 656 19054 732 19130
rect 656 18998 666 19054
rect 722 18998 732 19054
rect 656 18922 732 18998
rect 656 18866 666 18922
rect 722 18866 732 18922
rect 656 18790 732 18866
rect 656 18734 666 18790
rect 722 18734 732 18790
rect 656 18658 732 18734
rect 656 18602 666 18658
rect 722 18602 732 18658
rect 656 18526 732 18602
rect 656 18470 666 18526
rect 722 18470 732 18526
rect 656 18394 732 18470
rect 656 18338 666 18394
rect 722 18338 732 18394
rect 656 18262 732 18338
rect 656 18206 666 18262
rect 722 18206 732 18262
rect 656 18130 732 18206
rect 656 18074 666 18130
rect 722 18074 732 18130
rect 656 17998 732 18074
rect 656 17942 666 17998
rect 722 17942 732 17998
rect 656 17866 732 17942
rect 656 17810 666 17866
rect 722 17810 732 17866
rect 656 17734 732 17810
rect 656 17678 666 17734
rect 722 17678 732 17734
rect 656 17602 732 17678
rect 656 17546 666 17602
rect 722 17546 732 17602
rect 656 17470 732 17546
rect 656 17414 666 17470
rect 722 17414 732 17470
rect 656 16778 732 17414
rect 656 16722 666 16778
rect 722 16722 732 16778
rect 656 16646 732 16722
rect 656 16590 666 16646
rect 722 16590 732 16646
rect 656 16514 732 16590
rect 656 16458 666 16514
rect 722 16458 732 16514
rect 656 16382 732 16458
rect 656 16326 666 16382
rect 722 16326 732 16382
rect 656 16250 732 16326
rect 656 16194 666 16250
rect 722 16194 732 16250
rect 656 16118 732 16194
rect 656 16062 666 16118
rect 722 16062 732 16118
rect 656 15986 732 16062
rect 656 15930 666 15986
rect 722 15930 732 15986
rect 656 15854 732 15930
rect 656 15798 666 15854
rect 722 15798 732 15854
rect 656 15722 732 15798
rect 656 15666 666 15722
rect 722 15666 732 15722
rect 656 15590 732 15666
rect 656 15534 666 15590
rect 722 15534 732 15590
rect 656 15458 732 15534
rect 656 15402 666 15458
rect 722 15402 732 15458
rect 656 15326 732 15402
rect 656 15270 666 15326
rect 722 15270 732 15326
rect 656 15194 732 15270
rect 656 15138 666 15194
rect 722 15138 732 15194
rect 656 15062 732 15138
rect 656 15006 666 15062
rect 722 15006 732 15062
rect 656 14930 732 15006
rect 656 14874 666 14930
rect 722 14874 732 14930
rect 656 14798 732 14874
rect 656 14742 666 14798
rect 722 14742 732 14798
rect 656 14666 732 14742
rect 656 14610 666 14666
rect 722 14610 732 14666
rect 656 14534 732 14610
rect 656 14478 666 14534
rect 722 14478 732 14534
rect 656 14402 732 14478
rect 656 14346 666 14402
rect 722 14346 732 14402
rect 656 14270 732 14346
rect 656 14214 666 14270
rect 722 14214 732 14270
rect 656 14000 732 14214
rect 839 65000 915 69660
rect 839 64886 1000 65000
rect 839 64830 849 64886
rect 905 64830 1000 64886
rect 839 64762 1000 64830
rect 839 64706 849 64762
rect 905 64706 1000 64762
rect 839 64638 1000 64706
rect 839 64582 849 64638
rect 905 64582 1000 64638
rect 839 64514 1000 64582
rect 839 64458 849 64514
rect 905 64458 1000 64514
rect 839 64390 1000 64458
rect 839 64334 849 64390
rect 905 64334 1000 64390
rect 839 64266 1000 64334
rect 839 64210 849 64266
rect 905 64210 1000 64266
rect 839 64142 1000 64210
rect 839 64086 849 64142
rect 905 64086 1000 64142
rect 839 64018 1000 64086
rect 839 63962 849 64018
rect 905 63962 1000 64018
rect 839 63894 1000 63962
rect 839 63838 849 63894
rect 905 63838 1000 63894
rect 839 63770 1000 63838
rect 839 63714 849 63770
rect 905 63714 1000 63770
rect 839 63600 1000 63714
rect 839 50600 915 63600
rect 839 50486 1000 50600
rect 839 50430 849 50486
rect 905 50430 1000 50486
rect 839 50362 1000 50430
rect 839 50306 849 50362
rect 905 50306 1000 50362
rect 839 50238 1000 50306
rect 839 50182 849 50238
rect 905 50182 1000 50238
rect 839 50114 1000 50182
rect 839 50058 849 50114
rect 905 50058 1000 50114
rect 839 49990 1000 50058
rect 839 49934 849 49990
rect 905 49934 1000 49990
rect 839 49866 1000 49934
rect 839 49810 849 49866
rect 905 49810 1000 49866
rect 839 49742 1000 49810
rect 839 49686 849 49742
rect 905 49686 1000 49742
rect 839 49618 1000 49686
rect 839 49562 849 49618
rect 905 49562 1000 49618
rect 839 49494 1000 49562
rect 839 49438 849 49494
rect 905 49438 1000 49494
rect 839 49370 1000 49438
rect 839 49314 849 49370
rect 905 49314 1000 49370
rect 839 49200 1000 49314
rect 839 13494 915 49200
<< via2 >>
rect 666 69523 722 69579
rect 666 69391 722 69447
rect 666 69259 722 69315
rect 666 69127 722 69183
rect 666 68995 722 69051
rect 666 68863 722 68919
rect 666 68731 722 68787
rect 666 68599 722 68655
rect 666 68467 722 68523
rect 57 64884 113 64886
rect 57 64832 59 64884
rect 59 64832 111 64884
rect 111 64832 113 64884
rect 57 64830 113 64832
rect 57 64760 113 64762
rect 57 64708 59 64760
rect 59 64708 111 64760
rect 111 64708 113 64760
rect 57 64706 113 64708
rect 57 64636 113 64638
rect 57 64584 59 64636
rect 59 64584 111 64636
rect 111 64584 113 64636
rect 57 64582 113 64584
rect 57 64512 113 64514
rect 57 64460 59 64512
rect 59 64460 111 64512
rect 111 64460 113 64512
rect 57 64458 113 64460
rect 57 64388 113 64390
rect 57 64336 59 64388
rect 59 64336 111 64388
rect 111 64336 113 64388
rect 57 64334 113 64336
rect 57 64264 113 64266
rect 57 64212 59 64264
rect 59 64212 111 64264
rect 111 64212 113 64264
rect 57 64210 113 64212
rect 57 64140 113 64142
rect 57 64088 59 64140
rect 59 64088 111 64140
rect 111 64088 113 64140
rect 57 64086 113 64088
rect 57 64016 113 64018
rect 57 63964 59 64016
rect 59 63964 111 64016
rect 111 63964 113 64016
rect 57 63962 113 63964
rect 57 63892 113 63894
rect 57 63840 59 63892
rect 59 63840 111 63892
rect 111 63840 113 63892
rect 57 63838 113 63840
rect 57 63768 113 63770
rect 57 63716 59 63768
rect 59 63716 111 63768
rect 111 63716 113 63768
rect 57 63714 113 63716
rect 57 50484 113 50486
rect 57 50432 59 50484
rect 59 50432 111 50484
rect 111 50432 113 50484
rect 57 50430 113 50432
rect 57 50360 113 50362
rect 57 50308 59 50360
rect 59 50308 111 50360
rect 111 50308 113 50360
rect 57 50306 113 50308
rect 57 50236 113 50238
rect 57 50184 59 50236
rect 59 50184 111 50236
rect 111 50184 113 50236
rect 57 50182 113 50184
rect 57 50112 113 50114
rect 57 50060 59 50112
rect 59 50060 111 50112
rect 111 50060 113 50112
rect 57 50058 113 50060
rect 57 49988 113 49990
rect 57 49936 59 49988
rect 59 49936 111 49988
rect 111 49936 113 49988
rect 57 49934 113 49936
rect 57 49864 113 49866
rect 57 49812 59 49864
rect 59 49812 111 49864
rect 111 49812 113 49864
rect 57 49810 113 49812
rect 57 49740 113 49742
rect 57 49688 59 49740
rect 59 49688 111 49740
rect 111 49688 113 49740
rect 57 49686 113 49688
rect 57 49616 113 49618
rect 57 49564 59 49616
rect 59 49564 111 49616
rect 111 49564 113 49616
rect 57 49562 113 49564
rect 57 49492 113 49494
rect 57 49440 59 49492
rect 59 49440 111 49492
rect 111 49440 113 49492
rect 57 49438 113 49440
rect 57 49368 113 49370
rect 57 49316 59 49368
rect 59 49316 111 49368
rect 111 49316 113 49368
rect 57 49314 113 49316
rect 290 67994 346 68050
rect 290 67862 346 67918
rect 290 67730 346 67786
rect 290 67598 346 67654
rect 290 67466 346 67522
rect 290 67334 346 67390
rect 290 67202 346 67258
rect 290 67070 346 67126
rect 290 66938 346 66994
rect 666 66410 722 66466
rect 666 66278 722 66334
rect 666 66146 722 66202
rect 666 66014 722 66070
rect 666 65882 722 65938
rect 666 65750 722 65806
rect 666 65618 722 65674
rect 666 65486 722 65542
rect 666 65354 722 65410
rect 482 63197 538 63253
rect 482 63065 538 63121
rect 482 62933 538 62989
rect 482 62801 538 62857
rect 482 62669 538 62725
rect 482 62537 538 62593
rect 482 62405 538 62461
rect 482 62273 538 62329
rect 482 62141 538 62197
rect 290 60005 346 60061
rect 290 59873 346 59929
rect 290 59741 346 59797
rect 290 59609 346 59665
rect 290 59477 346 59533
rect 290 59345 346 59401
rect 290 59213 346 59269
rect 290 59081 346 59137
rect 290 58949 346 59005
rect 290 56823 346 56879
rect 290 56691 346 56747
rect 290 56559 346 56615
rect 290 56427 346 56483
rect 290 56295 346 56351
rect 290 56163 346 56219
rect 290 56031 346 56087
rect 290 55899 346 55955
rect 290 55767 346 55823
rect 290 55204 346 55260
rect 290 55072 346 55128
rect 290 54940 346 54996
rect 290 54808 346 54864
rect 290 54676 346 54732
rect 290 54544 346 54600
rect 290 54412 346 54468
rect 290 54280 346 54336
rect 290 54148 346 54204
rect 290 53613 346 53669
rect 290 53481 346 53537
rect 290 53349 346 53405
rect 290 53217 346 53273
rect 290 53085 346 53141
rect 290 52953 346 53009
rect 290 52821 346 52877
rect 290 52689 346 52745
rect 290 52557 346 52613
rect 666 61608 722 61664
rect 666 61476 722 61532
rect 666 61344 722 61400
rect 666 61212 722 61268
rect 666 61080 722 61136
rect 666 60948 722 61004
rect 666 60816 722 60872
rect 666 60684 722 60740
rect 666 60552 722 60608
rect 666 58397 722 58453
rect 666 58265 722 58321
rect 666 58133 722 58189
rect 666 58001 722 58057
rect 666 57869 722 57925
rect 666 57737 722 57793
rect 666 57605 722 57661
rect 666 57473 722 57529
rect 666 57341 722 57397
rect 482 52004 538 52060
rect 482 51872 538 51928
rect 482 51740 538 51796
rect 482 51608 538 51664
rect 482 51476 538 51532
rect 482 51344 538 51400
rect 482 51212 538 51268
rect 482 51080 538 51136
rect 482 50948 538 51004
rect 290 45537 346 45593
rect 290 45405 346 45461
rect 290 45273 346 45329
rect 290 45141 346 45197
rect 290 45009 346 45065
rect 290 44877 346 44933
rect 290 44745 346 44801
rect 290 44613 346 44669
rect 290 44481 346 44537
rect 290 44349 346 44405
rect 290 44217 346 44273
rect 290 44085 346 44141
rect 290 43953 346 44009
rect 290 43821 346 43877
rect 290 43689 346 43745
rect 290 43557 346 43613
rect 290 43425 346 43481
rect 290 43293 346 43349
rect 290 43161 346 43217
rect 290 43029 346 43085
rect 290 42395 346 42451
rect 290 42263 346 42319
rect 290 42131 346 42187
rect 290 41999 346 42055
rect 290 41867 346 41923
rect 290 41735 346 41791
rect 290 41603 346 41659
rect 290 41471 346 41527
rect 290 41339 346 41395
rect 290 39114 346 39170
rect 290 38982 346 39038
rect 290 38850 346 38906
rect 290 38718 346 38774
rect 290 38586 346 38642
rect 290 38454 346 38510
rect 290 38322 346 38378
rect 290 38190 346 38246
rect 290 38058 346 38114
rect 290 37926 346 37982
rect 290 37794 346 37850
rect 290 37662 346 37718
rect 290 37530 346 37586
rect 290 37398 346 37454
rect 290 37266 346 37322
rect 290 37134 346 37190
rect 290 37002 346 37058
rect 290 36870 346 36926
rect 290 36738 346 36794
rect 290 36606 346 36662
rect 290 35944 346 36000
rect 290 35812 346 35868
rect 290 35680 346 35736
rect 290 35548 346 35604
rect 290 35416 346 35472
rect 290 35284 346 35340
rect 290 35152 346 35208
rect 290 35020 346 35076
rect 290 34888 346 34944
rect 290 34756 346 34812
rect 290 34624 346 34680
rect 290 34492 346 34548
rect 290 34360 346 34416
rect 290 34228 346 34284
rect 290 34096 346 34152
rect 290 33964 346 34020
rect 290 33832 346 33888
rect 290 33700 346 33756
rect 290 33568 346 33624
rect 290 33436 346 33492
rect 290 32739 346 32795
rect 290 32607 346 32663
rect 290 32475 346 32531
rect 290 32343 346 32399
rect 290 32211 346 32267
rect 290 32079 346 32135
rect 290 31947 346 32003
rect 290 31815 346 31871
rect 290 31683 346 31739
rect 290 31551 346 31607
rect 290 31419 346 31475
rect 290 31287 346 31343
rect 290 31155 346 31211
rect 290 31023 346 31079
rect 290 30891 346 30947
rect 290 30759 346 30815
rect 290 30627 346 30683
rect 290 30495 346 30551
rect 290 30363 346 30419
rect 290 30231 346 30287
rect 290 29569 346 29625
rect 290 29437 346 29493
rect 290 29305 346 29361
rect 290 29173 346 29229
rect 290 29041 346 29097
rect 290 28909 346 28965
rect 290 28777 346 28833
rect 290 28645 346 28701
rect 290 28513 346 28569
rect 290 28381 346 28437
rect 290 28249 346 28305
rect 290 28117 346 28173
rect 290 27985 346 28041
rect 290 27853 346 27909
rect 290 27721 346 27777
rect 290 27589 346 27645
rect 290 27457 346 27513
rect 290 27325 346 27381
rect 290 27193 346 27249
rect 290 27061 346 27117
rect 290 24798 346 24854
rect 290 24666 346 24722
rect 290 24534 346 24590
rect 290 24402 346 24458
rect 290 24270 346 24326
rect 290 24138 346 24194
rect 290 24006 346 24062
rect 290 23874 346 23930
rect 290 23742 346 23798
rect 666 48754 722 48810
rect 666 48622 722 48678
rect 666 48490 722 48546
rect 666 48358 722 48414
rect 666 48226 722 48282
rect 666 48094 722 48150
rect 666 47962 722 48018
rect 666 47830 722 47886
rect 666 47698 722 47754
rect 666 47566 722 47622
rect 666 47434 722 47490
rect 666 47302 722 47358
rect 666 47170 722 47226
rect 666 47038 722 47094
rect 666 46906 722 46962
rect 666 46774 722 46830
rect 666 46642 722 46698
rect 666 46510 722 46566
rect 666 46378 722 46434
rect 666 46246 722 46302
rect 666 40827 722 40883
rect 666 40695 722 40751
rect 666 40563 722 40619
rect 666 40431 722 40487
rect 666 40299 722 40355
rect 666 40167 722 40223
rect 666 40035 722 40091
rect 666 39903 722 39959
rect 666 39771 722 39827
rect 666 26429 722 26485
rect 666 26297 722 26353
rect 666 26165 722 26221
rect 666 26033 722 26089
rect 666 25901 722 25957
rect 666 25769 722 25825
rect 666 25637 722 25693
rect 666 25505 722 25561
rect 666 25373 722 25429
rect 666 23134 722 23190
rect 666 23002 722 23058
rect 666 22870 722 22926
rect 666 22738 722 22794
rect 666 22606 722 22662
rect 666 22474 722 22530
rect 666 22342 722 22398
rect 666 22210 722 22266
rect 666 22078 722 22134
rect 666 21946 722 22002
rect 666 21814 722 21870
rect 666 21682 722 21738
rect 666 21550 722 21606
rect 666 21418 722 21474
rect 666 21286 722 21342
rect 666 21154 722 21210
rect 666 21022 722 21078
rect 666 20890 722 20946
rect 666 20758 722 20814
rect 666 20626 722 20682
rect 666 19922 722 19978
rect 666 19790 722 19846
rect 666 19658 722 19714
rect 666 19526 722 19582
rect 666 19394 722 19450
rect 666 19262 722 19318
rect 666 19130 722 19186
rect 666 18998 722 19054
rect 666 18866 722 18922
rect 666 18734 722 18790
rect 666 18602 722 18658
rect 666 18470 722 18526
rect 666 18338 722 18394
rect 666 18206 722 18262
rect 666 18074 722 18130
rect 666 17942 722 17998
rect 666 17810 722 17866
rect 666 17678 722 17734
rect 666 17546 722 17602
rect 666 17414 722 17470
rect 666 16722 722 16778
rect 666 16590 722 16646
rect 666 16458 722 16514
rect 666 16326 722 16382
rect 666 16194 722 16250
rect 666 16062 722 16118
rect 666 15930 722 15986
rect 666 15798 722 15854
rect 666 15666 722 15722
rect 666 15534 722 15590
rect 666 15402 722 15458
rect 666 15270 722 15326
rect 666 15138 722 15194
rect 666 15006 722 15062
rect 666 14874 722 14930
rect 666 14742 722 14798
rect 666 14610 722 14666
rect 666 14478 722 14534
rect 666 14346 722 14402
rect 666 14214 722 14270
rect 849 64884 905 64886
rect 849 64832 851 64884
rect 851 64832 903 64884
rect 903 64832 905 64884
rect 849 64830 905 64832
rect 849 64760 905 64762
rect 849 64708 851 64760
rect 851 64708 903 64760
rect 903 64708 905 64760
rect 849 64706 905 64708
rect 849 64636 905 64638
rect 849 64584 851 64636
rect 851 64584 903 64636
rect 903 64584 905 64636
rect 849 64582 905 64584
rect 849 64512 905 64514
rect 849 64460 851 64512
rect 851 64460 903 64512
rect 903 64460 905 64512
rect 849 64458 905 64460
rect 849 64388 905 64390
rect 849 64336 851 64388
rect 851 64336 903 64388
rect 903 64336 905 64388
rect 849 64334 905 64336
rect 849 64264 905 64266
rect 849 64212 851 64264
rect 851 64212 903 64264
rect 903 64212 905 64264
rect 849 64210 905 64212
rect 849 64140 905 64142
rect 849 64088 851 64140
rect 851 64088 903 64140
rect 903 64088 905 64140
rect 849 64086 905 64088
rect 849 64016 905 64018
rect 849 63964 851 64016
rect 851 63964 903 64016
rect 903 63964 905 64016
rect 849 63962 905 63964
rect 849 63892 905 63894
rect 849 63840 851 63892
rect 851 63840 903 63892
rect 903 63840 905 63892
rect 849 63838 905 63840
rect 849 63768 905 63770
rect 849 63716 851 63768
rect 851 63716 903 63768
rect 903 63716 905 63768
rect 849 63714 905 63716
rect 849 50484 905 50486
rect 849 50432 851 50484
rect 851 50432 903 50484
rect 903 50432 905 50484
rect 849 50430 905 50432
rect 849 50360 905 50362
rect 849 50308 851 50360
rect 851 50308 903 50360
rect 903 50308 905 50360
rect 849 50306 905 50308
rect 849 50236 905 50238
rect 849 50184 851 50236
rect 851 50184 903 50236
rect 903 50184 905 50236
rect 849 50182 905 50184
rect 849 50112 905 50114
rect 849 50060 851 50112
rect 851 50060 903 50112
rect 903 50060 905 50112
rect 849 50058 905 50060
rect 849 49988 905 49990
rect 849 49936 851 49988
rect 851 49936 903 49988
rect 903 49936 905 49988
rect 849 49934 905 49936
rect 849 49864 905 49866
rect 849 49812 851 49864
rect 851 49812 903 49864
rect 903 49812 905 49864
rect 849 49810 905 49812
rect 849 49740 905 49742
rect 849 49688 851 49740
rect 851 49688 903 49740
rect 903 49688 905 49740
rect 849 49686 905 49688
rect 849 49616 905 49618
rect 849 49564 851 49616
rect 851 49564 903 49616
rect 903 49564 905 49616
rect 849 49562 905 49564
rect 849 49492 905 49494
rect 849 49440 851 49492
rect 851 49440 903 49492
rect 903 49440 905 49492
rect 849 49438 905 49440
rect 849 49368 905 49370
rect 849 49316 851 49368
rect 851 49316 903 49368
rect 903 49316 905 49368
rect 849 49314 905 49316
<< metal3 >>
rect 0 69579 1000 69678
rect 0 69523 666 69579
rect 722 69523 1000 69579
rect 0 69447 1000 69523
rect 0 69391 666 69447
rect 722 69391 1000 69447
rect 0 69315 1000 69391
rect 0 69259 666 69315
rect 722 69259 1000 69315
rect 0 69183 1000 69259
rect 0 69127 666 69183
rect 722 69127 1000 69183
rect 0 69051 1000 69127
rect 0 68995 666 69051
rect 722 68995 1000 69051
rect 0 68919 1000 68995
rect 0 68863 666 68919
rect 722 68863 1000 68919
rect 0 68787 1000 68863
rect 0 68731 666 68787
rect 722 68731 1000 68787
rect 0 68655 1000 68731
rect 0 68599 666 68655
rect 722 68599 1000 68655
rect 0 68523 1000 68599
rect 0 68467 666 68523
rect 722 68467 1000 68523
rect 0 68400 1000 68467
rect 0 68050 1000 68200
rect 0 67994 290 68050
rect 346 67994 1000 68050
rect 0 67918 1000 67994
rect 0 67862 290 67918
rect 346 67862 1000 67918
rect 0 67786 1000 67862
rect 0 67730 290 67786
rect 346 67730 1000 67786
rect 0 67654 1000 67730
rect 0 67598 290 67654
rect 346 67598 1000 67654
rect 0 67522 1000 67598
rect 0 67466 290 67522
rect 346 67466 1000 67522
rect 0 67390 1000 67466
rect 0 67334 290 67390
rect 346 67334 1000 67390
rect 0 67258 1000 67334
rect 0 67202 290 67258
rect 346 67202 1000 67258
rect 0 67126 1000 67202
rect 0 67070 290 67126
rect 346 67070 1000 67126
rect 0 66994 1000 67070
rect 0 66938 290 66994
rect 346 66938 1000 66994
rect 0 66800 1000 66938
rect 0 66466 1000 66600
rect 0 66410 666 66466
rect 722 66410 1000 66466
rect 0 66334 1000 66410
rect 0 66278 666 66334
rect 722 66278 1000 66334
rect 0 66202 1000 66278
rect 0 66146 666 66202
rect 722 66146 1000 66202
rect 0 66070 1000 66146
rect 0 66014 666 66070
rect 722 66014 1000 66070
rect 0 65938 1000 66014
rect 0 65882 666 65938
rect 722 65882 1000 65938
rect 0 65806 1000 65882
rect 0 65750 666 65806
rect 722 65750 1000 65806
rect 0 65674 1000 65750
rect 0 65618 666 65674
rect 722 65618 1000 65674
rect 0 65542 1000 65618
rect 0 65486 666 65542
rect 722 65486 1000 65542
rect 0 65410 1000 65486
rect 0 65354 666 65410
rect 722 65354 1000 65410
rect 0 65200 1000 65354
rect 0 64886 1000 65000
rect 0 64830 57 64886
rect 113 64830 849 64886
rect 905 64830 1000 64886
rect 0 64762 1000 64830
rect 0 64706 57 64762
rect 113 64706 849 64762
rect 905 64706 1000 64762
rect 0 64638 1000 64706
rect 0 64582 57 64638
rect 113 64582 849 64638
rect 905 64582 1000 64638
rect 0 64514 1000 64582
rect 0 64458 57 64514
rect 113 64458 849 64514
rect 905 64458 1000 64514
rect 0 64390 1000 64458
rect 0 64334 57 64390
rect 113 64334 849 64390
rect 905 64334 1000 64390
rect 0 64266 1000 64334
rect 0 64210 57 64266
rect 113 64210 849 64266
rect 905 64210 1000 64266
rect 0 64142 1000 64210
rect 0 64086 57 64142
rect 113 64086 849 64142
rect 905 64086 1000 64142
rect 0 64018 1000 64086
rect 0 63962 57 64018
rect 113 63962 849 64018
rect 905 63962 1000 64018
rect 0 63894 1000 63962
rect 0 63838 57 63894
rect 113 63838 849 63894
rect 905 63838 1000 63894
rect 0 63770 1000 63838
rect 0 63714 57 63770
rect 113 63714 849 63770
rect 905 63714 1000 63770
rect 0 63600 1000 63714
rect 0 63253 1000 63400
rect 0 63197 482 63253
rect 538 63197 1000 63253
rect 0 63121 1000 63197
rect 0 63065 482 63121
rect 538 63065 1000 63121
rect 0 62989 1000 63065
rect 0 62933 482 62989
rect 538 62933 1000 62989
rect 0 62857 1000 62933
rect 0 62801 482 62857
rect 538 62801 1000 62857
rect 0 62725 1000 62801
rect 0 62669 482 62725
rect 538 62669 1000 62725
rect 0 62593 1000 62669
rect 0 62537 482 62593
rect 538 62537 1000 62593
rect 0 62461 1000 62537
rect 0 62405 482 62461
rect 538 62405 1000 62461
rect 0 62329 1000 62405
rect 0 62273 482 62329
rect 538 62273 1000 62329
rect 0 62197 1000 62273
rect 0 62141 482 62197
rect 538 62141 1000 62197
rect 0 62000 1000 62141
rect 0 61664 1000 61800
rect 0 61608 666 61664
rect 722 61608 1000 61664
rect 0 61532 1000 61608
rect 0 61476 666 61532
rect 722 61476 1000 61532
rect 0 61400 1000 61476
rect 0 61344 666 61400
rect 722 61344 1000 61400
rect 0 61268 1000 61344
rect 0 61212 666 61268
rect 722 61212 1000 61268
rect 0 61136 1000 61212
rect 0 61080 666 61136
rect 722 61080 1000 61136
rect 0 61004 1000 61080
rect 0 60948 666 61004
rect 722 60948 1000 61004
rect 0 60872 1000 60948
rect 0 60816 666 60872
rect 722 60816 1000 60872
rect 0 60740 1000 60816
rect 0 60684 666 60740
rect 722 60684 1000 60740
rect 0 60608 1000 60684
rect 0 60552 666 60608
rect 722 60552 1000 60608
rect 0 60400 1000 60552
rect 0 60061 1000 60200
rect 0 60005 290 60061
rect 346 60005 1000 60061
rect 0 59929 1000 60005
rect 0 59873 290 59929
rect 346 59873 1000 59929
rect 0 59797 1000 59873
rect 0 59741 290 59797
rect 346 59741 1000 59797
rect 0 59665 1000 59741
rect 0 59609 290 59665
rect 346 59609 1000 59665
rect 0 59533 1000 59609
rect 0 59477 290 59533
rect 346 59477 1000 59533
rect 0 59401 1000 59477
rect 0 59345 290 59401
rect 346 59345 1000 59401
rect 0 59269 1000 59345
rect 0 59213 290 59269
rect 346 59213 1000 59269
rect 0 59137 1000 59213
rect 0 59081 290 59137
rect 346 59081 1000 59137
rect 0 59005 1000 59081
rect 0 58949 290 59005
rect 346 58949 1000 59005
rect 0 58800 1000 58949
rect 0 58453 1000 58600
rect 0 58397 666 58453
rect 722 58397 1000 58453
rect 0 58321 1000 58397
rect 0 58265 666 58321
rect 722 58265 1000 58321
rect 0 58189 1000 58265
rect 0 58133 666 58189
rect 722 58133 1000 58189
rect 0 58057 1000 58133
rect 0 58001 666 58057
rect 722 58001 1000 58057
rect 0 57925 1000 58001
rect 0 57869 666 57925
rect 722 57869 1000 57925
rect 0 57793 1000 57869
rect 0 57737 666 57793
rect 722 57737 1000 57793
rect 0 57661 1000 57737
rect 0 57605 666 57661
rect 722 57605 1000 57661
rect 0 57529 1000 57605
rect 0 57473 666 57529
rect 722 57473 1000 57529
rect 0 57397 1000 57473
rect 0 57341 666 57397
rect 722 57341 1000 57397
rect 0 57200 1000 57341
rect 0 56879 1000 57000
rect 0 56823 290 56879
rect 346 56823 1000 56879
rect 0 56747 1000 56823
rect 0 56691 290 56747
rect 346 56691 1000 56747
rect 0 56615 1000 56691
rect 0 56559 290 56615
rect 346 56559 1000 56615
rect 0 56483 1000 56559
rect 0 56427 290 56483
rect 346 56427 1000 56483
rect 0 56351 1000 56427
rect 0 56295 290 56351
rect 346 56295 1000 56351
rect 0 56219 1000 56295
rect 0 56163 290 56219
rect 346 56163 1000 56219
rect 0 56087 1000 56163
rect 0 56031 290 56087
rect 346 56031 1000 56087
rect 0 55955 1000 56031
rect 0 55899 290 55955
rect 346 55899 1000 55955
rect 0 55823 1000 55899
rect 0 55767 290 55823
rect 346 55767 1000 55823
rect 0 55600 1000 55767
rect 0 55260 1000 55400
rect 0 55204 290 55260
rect 346 55204 1000 55260
rect 0 55128 1000 55204
rect 0 55072 290 55128
rect 346 55072 1000 55128
rect 0 54996 1000 55072
rect 0 54940 290 54996
rect 346 54940 1000 54996
rect 0 54864 1000 54940
rect 0 54808 290 54864
rect 346 54808 1000 54864
rect 0 54732 1000 54808
rect 0 54676 290 54732
rect 346 54676 1000 54732
rect 0 54600 1000 54676
rect 0 54544 290 54600
rect 346 54544 1000 54600
rect 0 54468 1000 54544
rect 0 54412 290 54468
rect 346 54412 1000 54468
rect 0 54336 1000 54412
rect 0 54280 290 54336
rect 346 54280 1000 54336
rect 0 54204 1000 54280
rect 0 54148 290 54204
rect 346 54148 1000 54204
rect 0 54000 1000 54148
rect 0 53669 1000 53800
rect 0 53613 290 53669
rect 346 53613 1000 53669
rect 0 53537 1000 53613
rect 0 53481 290 53537
rect 346 53481 1000 53537
rect 0 53405 1000 53481
rect 0 53349 290 53405
rect 346 53349 1000 53405
rect 0 53273 1000 53349
rect 0 53217 290 53273
rect 346 53217 1000 53273
rect 0 53141 1000 53217
rect 0 53085 290 53141
rect 346 53085 1000 53141
rect 0 53009 1000 53085
rect 0 52953 290 53009
rect 346 52953 1000 53009
rect 0 52877 1000 52953
rect 0 52821 290 52877
rect 346 52821 1000 52877
rect 0 52745 1000 52821
rect 0 52689 290 52745
rect 346 52689 1000 52745
rect 0 52613 1000 52689
rect 0 52557 290 52613
rect 346 52557 1000 52613
rect 0 52400 1000 52557
rect 0 52060 1000 52200
rect 0 52004 482 52060
rect 538 52004 1000 52060
rect 0 51928 1000 52004
rect 0 51872 482 51928
rect 538 51872 1000 51928
rect 0 51796 1000 51872
rect 0 51740 482 51796
rect 538 51740 1000 51796
rect 0 51664 1000 51740
rect 0 51608 482 51664
rect 538 51608 1000 51664
rect 0 51532 1000 51608
rect 0 51476 482 51532
rect 538 51476 1000 51532
rect 0 51400 1000 51476
rect 0 51344 482 51400
rect 538 51344 1000 51400
rect 0 51268 1000 51344
rect 0 51212 482 51268
rect 538 51212 1000 51268
rect 0 51136 1000 51212
rect 0 51080 482 51136
rect 538 51080 1000 51136
rect 0 51004 1000 51080
rect 0 50948 482 51004
rect 538 50948 1000 51004
rect 0 50800 1000 50948
rect 0 50486 1000 50600
rect 0 50430 57 50486
rect 113 50430 849 50486
rect 905 50430 1000 50486
rect 0 50362 1000 50430
rect 0 50306 57 50362
rect 113 50306 849 50362
rect 905 50306 1000 50362
rect 0 50238 1000 50306
rect 0 50182 57 50238
rect 113 50182 849 50238
rect 905 50182 1000 50238
rect 0 50114 1000 50182
rect 0 50058 57 50114
rect 113 50058 849 50114
rect 905 50058 1000 50114
rect 0 49990 1000 50058
rect 0 49934 57 49990
rect 113 49934 849 49990
rect 905 49934 1000 49990
rect 0 49866 1000 49934
rect 0 49810 57 49866
rect 113 49810 849 49866
rect 905 49810 1000 49866
rect 0 49742 1000 49810
rect 0 49686 57 49742
rect 113 49686 849 49742
rect 905 49686 1000 49742
rect 0 49618 1000 49686
rect 0 49562 57 49618
rect 113 49562 849 49618
rect 905 49562 1000 49618
rect 0 49494 1000 49562
rect 0 49438 57 49494
rect 113 49438 849 49494
rect 905 49438 1000 49494
rect 0 49370 1000 49438
rect 0 49314 57 49370
rect 113 49314 849 49370
rect 905 49314 1000 49370
rect 0 49200 1000 49314
rect 0 48810 1000 49000
rect 0 48754 666 48810
rect 722 48754 1000 48810
rect 0 48678 1000 48754
rect 0 48622 666 48678
rect 722 48622 1000 48678
rect 0 48546 1000 48622
rect 0 48490 666 48546
rect 722 48490 1000 48546
rect 0 48414 1000 48490
rect 0 48358 666 48414
rect 722 48358 1000 48414
rect 0 48282 1000 48358
rect 0 48226 666 48282
rect 722 48226 1000 48282
rect 0 48150 1000 48226
rect 0 48094 666 48150
rect 722 48094 1000 48150
rect 0 48018 1000 48094
rect 0 47962 666 48018
rect 722 47962 1000 48018
rect 0 47886 1000 47962
rect 0 47830 666 47886
rect 722 47830 1000 47886
rect 0 47754 1000 47830
rect 0 47698 666 47754
rect 722 47698 1000 47754
rect 0 47622 1000 47698
rect 0 47566 666 47622
rect 722 47566 1000 47622
rect 0 47490 1000 47566
rect 0 47434 666 47490
rect 722 47434 1000 47490
rect 0 47358 1000 47434
rect 0 47302 666 47358
rect 722 47302 1000 47358
rect 0 47226 1000 47302
rect 0 47170 666 47226
rect 722 47170 1000 47226
rect 0 47094 1000 47170
rect 0 47038 666 47094
rect 722 47038 1000 47094
rect 0 46962 1000 47038
rect 0 46906 666 46962
rect 722 46906 1000 46962
rect 0 46830 1000 46906
rect 0 46774 666 46830
rect 722 46774 1000 46830
rect 0 46698 1000 46774
rect 0 46642 666 46698
rect 722 46642 1000 46698
rect 0 46566 1000 46642
rect 0 46510 666 46566
rect 722 46510 1000 46566
rect 0 46434 1000 46510
rect 0 46378 666 46434
rect 722 46378 1000 46434
rect 0 46302 1000 46378
rect 0 46246 666 46302
rect 722 46246 1000 46302
rect 0 46000 1000 46246
rect 0 45593 1000 45800
rect 0 45537 290 45593
rect 346 45537 1000 45593
rect 0 45461 1000 45537
rect 0 45405 290 45461
rect 346 45405 1000 45461
rect 0 45329 1000 45405
rect 0 45273 290 45329
rect 346 45273 1000 45329
rect 0 45197 1000 45273
rect 0 45141 290 45197
rect 346 45141 1000 45197
rect 0 45065 1000 45141
rect 0 45009 290 45065
rect 346 45009 1000 45065
rect 0 44933 1000 45009
rect 0 44877 290 44933
rect 346 44877 1000 44933
rect 0 44801 1000 44877
rect 0 44745 290 44801
rect 346 44745 1000 44801
rect 0 44669 1000 44745
rect 0 44613 290 44669
rect 346 44613 1000 44669
rect 0 44537 1000 44613
rect 0 44481 290 44537
rect 346 44481 1000 44537
rect 0 44405 1000 44481
rect 0 44349 290 44405
rect 346 44349 1000 44405
rect 0 44273 1000 44349
rect 0 44217 290 44273
rect 346 44217 1000 44273
rect 0 44141 1000 44217
rect 0 44085 290 44141
rect 346 44085 1000 44141
rect 0 44009 1000 44085
rect 0 43953 290 44009
rect 346 43953 1000 44009
rect 0 43877 1000 43953
rect 0 43821 290 43877
rect 346 43821 1000 43877
rect 0 43745 1000 43821
rect 0 43689 290 43745
rect 346 43689 1000 43745
rect 0 43613 1000 43689
rect 0 43557 290 43613
rect 346 43557 1000 43613
rect 0 43481 1000 43557
rect 0 43425 290 43481
rect 346 43425 1000 43481
rect 0 43349 1000 43425
rect 0 43293 290 43349
rect 346 43293 1000 43349
rect 0 43217 1000 43293
rect 0 43161 290 43217
rect 346 43161 1000 43217
rect 0 43085 1000 43161
rect 0 43029 290 43085
rect 346 43029 1000 43085
rect 0 42800 1000 43029
rect 0 42451 1000 42600
rect 0 42395 290 42451
rect 346 42395 1000 42451
rect 0 42319 1000 42395
rect 0 42263 290 42319
rect 346 42263 1000 42319
rect 0 42187 1000 42263
rect 0 42131 290 42187
rect 346 42131 1000 42187
rect 0 42055 1000 42131
rect 0 41999 290 42055
rect 346 41999 1000 42055
rect 0 41923 1000 41999
rect 0 41867 290 41923
rect 346 41867 1000 41923
rect 0 41791 1000 41867
rect 0 41735 290 41791
rect 346 41735 1000 41791
rect 0 41659 1000 41735
rect 0 41603 290 41659
rect 346 41603 1000 41659
rect 0 41527 1000 41603
rect 0 41471 290 41527
rect 346 41471 1000 41527
rect 0 41395 1000 41471
rect 0 41339 290 41395
rect 346 41339 1000 41395
rect 0 41200 1000 41339
rect 0 40883 1000 41000
rect 0 40827 666 40883
rect 722 40827 1000 40883
rect 0 40751 1000 40827
rect 0 40695 666 40751
rect 722 40695 1000 40751
rect 0 40619 1000 40695
rect 0 40563 666 40619
rect 722 40563 1000 40619
rect 0 40487 1000 40563
rect 0 40431 666 40487
rect 722 40431 1000 40487
rect 0 40355 1000 40431
rect 0 40299 666 40355
rect 722 40299 1000 40355
rect 0 40223 1000 40299
rect 0 40167 666 40223
rect 722 40167 1000 40223
rect 0 40091 1000 40167
rect 0 40035 666 40091
rect 722 40035 1000 40091
rect 0 39959 1000 40035
rect 0 39903 666 39959
rect 722 39903 1000 39959
rect 0 39827 1000 39903
rect 0 39771 666 39827
rect 722 39771 1000 39827
rect 0 39600 1000 39771
rect 0 39170 1000 39400
rect 0 39114 290 39170
rect 346 39114 1000 39170
rect 0 39038 1000 39114
rect 0 38982 290 39038
rect 346 38982 1000 39038
rect 0 38906 1000 38982
rect 0 38850 290 38906
rect 346 38850 1000 38906
rect 0 38774 1000 38850
rect 0 38718 290 38774
rect 346 38718 1000 38774
rect 0 38642 1000 38718
rect 0 38586 290 38642
rect 346 38586 1000 38642
rect 0 38510 1000 38586
rect 0 38454 290 38510
rect 346 38454 1000 38510
rect 0 38378 1000 38454
rect 0 38322 290 38378
rect 346 38322 1000 38378
rect 0 38246 1000 38322
rect 0 38190 290 38246
rect 346 38190 1000 38246
rect 0 38114 1000 38190
rect 0 38058 290 38114
rect 346 38058 1000 38114
rect 0 37982 1000 38058
rect 0 37926 290 37982
rect 346 37926 1000 37982
rect 0 37850 1000 37926
rect 0 37794 290 37850
rect 346 37794 1000 37850
rect 0 37718 1000 37794
rect 0 37662 290 37718
rect 346 37662 1000 37718
rect 0 37586 1000 37662
rect 0 37530 290 37586
rect 346 37530 1000 37586
rect 0 37454 1000 37530
rect 0 37398 290 37454
rect 346 37398 1000 37454
rect 0 37322 1000 37398
rect 0 37266 290 37322
rect 346 37266 1000 37322
rect 0 37190 1000 37266
rect 0 37134 290 37190
rect 346 37134 1000 37190
rect 0 37058 1000 37134
rect 0 37002 290 37058
rect 346 37002 1000 37058
rect 0 36926 1000 37002
rect 0 36870 290 36926
rect 346 36870 1000 36926
rect 0 36794 1000 36870
rect 0 36738 290 36794
rect 346 36738 1000 36794
rect 0 36662 1000 36738
rect 0 36606 290 36662
rect 346 36606 1000 36662
rect 0 36400 1000 36606
rect 0 36000 1000 36200
rect 0 35944 290 36000
rect 346 35944 1000 36000
rect 0 35868 1000 35944
rect 0 35812 290 35868
rect 346 35812 1000 35868
rect 0 35736 1000 35812
rect 0 35680 290 35736
rect 346 35680 1000 35736
rect 0 35604 1000 35680
rect 0 35548 290 35604
rect 346 35548 1000 35604
rect 0 35472 1000 35548
rect 0 35416 290 35472
rect 346 35416 1000 35472
rect 0 35340 1000 35416
rect 0 35284 290 35340
rect 346 35284 1000 35340
rect 0 35208 1000 35284
rect 0 35152 290 35208
rect 346 35152 1000 35208
rect 0 35076 1000 35152
rect 0 35020 290 35076
rect 346 35020 1000 35076
rect 0 34944 1000 35020
rect 0 34888 290 34944
rect 346 34888 1000 34944
rect 0 34812 1000 34888
rect 0 34756 290 34812
rect 346 34756 1000 34812
rect 0 34680 1000 34756
rect 0 34624 290 34680
rect 346 34624 1000 34680
rect 0 34548 1000 34624
rect 0 34492 290 34548
rect 346 34492 1000 34548
rect 0 34416 1000 34492
rect 0 34360 290 34416
rect 346 34360 1000 34416
rect 0 34284 1000 34360
rect 0 34228 290 34284
rect 346 34228 1000 34284
rect 0 34152 1000 34228
rect 0 34096 290 34152
rect 346 34096 1000 34152
rect 0 34020 1000 34096
rect 0 33964 290 34020
rect 346 33964 1000 34020
rect 0 33888 1000 33964
rect 0 33832 290 33888
rect 346 33832 1000 33888
rect 0 33756 1000 33832
rect 0 33700 290 33756
rect 346 33700 1000 33756
rect 0 33624 1000 33700
rect 0 33568 290 33624
rect 346 33568 1000 33624
rect 0 33492 1000 33568
rect 0 33436 290 33492
rect 346 33436 1000 33492
rect 0 33200 1000 33436
rect 0 32795 1000 33000
rect 0 32739 290 32795
rect 346 32739 1000 32795
rect 0 32663 1000 32739
rect 0 32607 290 32663
rect 346 32607 1000 32663
rect 0 32531 1000 32607
rect 0 32475 290 32531
rect 346 32475 1000 32531
rect 0 32399 1000 32475
rect 0 32343 290 32399
rect 346 32343 1000 32399
rect 0 32267 1000 32343
rect 0 32211 290 32267
rect 346 32211 1000 32267
rect 0 32135 1000 32211
rect 0 32079 290 32135
rect 346 32079 1000 32135
rect 0 32003 1000 32079
rect 0 31947 290 32003
rect 346 31947 1000 32003
rect 0 31871 1000 31947
rect 0 31815 290 31871
rect 346 31815 1000 31871
rect 0 31739 1000 31815
rect 0 31683 290 31739
rect 346 31683 1000 31739
rect 0 31607 1000 31683
rect 0 31551 290 31607
rect 346 31551 1000 31607
rect 0 31475 1000 31551
rect 0 31419 290 31475
rect 346 31419 1000 31475
rect 0 31343 1000 31419
rect 0 31287 290 31343
rect 346 31287 1000 31343
rect 0 31211 1000 31287
rect 0 31155 290 31211
rect 346 31155 1000 31211
rect 0 31079 1000 31155
rect 0 31023 290 31079
rect 346 31023 1000 31079
rect 0 30947 1000 31023
rect 0 30891 290 30947
rect 346 30891 1000 30947
rect 0 30815 1000 30891
rect 0 30759 290 30815
rect 346 30759 1000 30815
rect 0 30683 1000 30759
rect 0 30627 290 30683
rect 346 30627 1000 30683
rect 0 30551 1000 30627
rect 0 30495 290 30551
rect 346 30495 1000 30551
rect 0 30419 1000 30495
rect 0 30363 290 30419
rect 346 30363 1000 30419
rect 0 30287 1000 30363
rect 0 30231 290 30287
rect 346 30231 1000 30287
rect 0 30000 1000 30231
rect 0 29625 1000 29800
rect 0 29569 290 29625
rect 346 29569 1000 29625
rect 0 29493 1000 29569
rect 0 29437 290 29493
rect 346 29437 1000 29493
rect 0 29361 1000 29437
rect 0 29305 290 29361
rect 346 29305 1000 29361
rect 0 29229 1000 29305
rect 0 29173 290 29229
rect 346 29173 1000 29229
rect 0 29097 1000 29173
rect 0 29041 290 29097
rect 346 29041 1000 29097
rect 0 28965 1000 29041
rect 0 28909 290 28965
rect 346 28909 1000 28965
rect 0 28833 1000 28909
rect 0 28777 290 28833
rect 346 28777 1000 28833
rect 0 28701 1000 28777
rect 0 28645 290 28701
rect 346 28645 1000 28701
rect 0 28569 1000 28645
rect 0 28513 290 28569
rect 346 28513 1000 28569
rect 0 28437 1000 28513
rect 0 28381 290 28437
rect 346 28381 1000 28437
rect 0 28305 1000 28381
rect 0 28249 290 28305
rect 346 28249 1000 28305
rect 0 28173 1000 28249
rect 0 28117 290 28173
rect 346 28117 1000 28173
rect 0 28041 1000 28117
rect 0 27985 290 28041
rect 346 27985 1000 28041
rect 0 27909 1000 27985
rect 0 27853 290 27909
rect 346 27853 1000 27909
rect 0 27777 1000 27853
rect 0 27721 290 27777
rect 346 27721 1000 27777
rect 0 27645 1000 27721
rect 0 27589 290 27645
rect 346 27589 1000 27645
rect 0 27513 1000 27589
rect 0 27457 290 27513
rect 346 27457 1000 27513
rect 0 27381 1000 27457
rect 0 27325 290 27381
rect 346 27325 1000 27381
rect 0 27249 1000 27325
rect 0 27193 290 27249
rect 346 27193 1000 27249
rect 0 27117 1000 27193
rect 0 27061 290 27117
rect 346 27061 1000 27117
rect 0 26800 1000 27061
rect 0 26485 1000 26600
rect 0 26429 666 26485
rect 722 26429 1000 26485
rect 0 26353 1000 26429
rect 0 26297 666 26353
rect 722 26297 1000 26353
rect 0 26221 1000 26297
rect 0 26165 666 26221
rect 722 26165 1000 26221
rect 0 26089 1000 26165
rect 0 26033 666 26089
rect 722 26033 1000 26089
rect 0 25957 1000 26033
rect 0 25901 666 25957
rect 722 25901 1000 25957
rect 0 25825 1000 25901
rect 0 25769 666 25825
rect 722 25769 1000 25825
rect 0 25693 1000 25769
rect 0 25637 666 25693
rect 722 25637 1000 25693
rect 0 25561 1000 25637
rect 0 25505 666 25561
rect 722 25505 1000 25561
rect 0 25429 1000 25505
rect 0 25373 666 25429
rect 722 25373 1000 25429
rect 0 25200 1000 25373
rect 0 24854 1000 25000
rect 0 24798 290 24854
rect 346 24798 1000 24854
rect 0 24722 1000 24798
rect 0 24666 290 24722
rect 346 24666 1000 24722
rect 0 24590 1000 24666
rect 0 24534 290 24590
rect 346 24534 1000 24590
rect 0 24458 1000 24534
rect 0 24402 290 24458
rect 346 24402 1000 24458
rect 0 24326 1000 24402
rect 0 24270 290 24326
rect 346 24270 1000 24326
rect 0 24194 1000 24270
rect 0 24138 290 24194
rect 346 24138 1000 24194
rect 0 24062 1000 24138
rect 0 24006 290 24062
rect 346 24006 1000 24062
rect 0 23930 1000 24006
rect 0 23874 290 23930
rect 346 23874 1000 23930
rect 0 23798 1000 23874
rect 0 23742 290 23798
rect 346 23742 1000 23798
rect 0 23600 1000 23742
rect 0 23190 1000 23400
rect 0 23134 666 23190
rect 722 23134 1000 23190
rect 0 23058 1000 23134
rect 0 23002 666 23058
rect 722 23002 1000 23058
rect 0 22926 1000 23002
rect 0 22870 666 22926
rect 722 22870 1000 22926
rect 0 22794 1000 22870
rect 0 22738 666 22794
rect 722 22738 1000 22794
rect 0 22662 1000 22738
rect 0 22606 666 22662
rect 722 22606 1000 22662
rect 0 22530 1000 22606
rect 0 22474 666 22530
rect 722 22474 1000 22530
rect 0 22398 1000 22474
rect 0 22342 666 22398
rect 722 22342 1000 22398
rect 0 22266 1000 22342
rect 0 22210 666 22266
rect 722 22210 1000 22266
rect 0 22134 1000 22210
rect 0 22078 666 22134
rect 722 22078 1000 22134
rect 0 22002 1000 22078
rect 0 21946 666 22002
rect 722 21946 1000 22002
rect 0 21870 1000 21946
rect 0 21814 666 21870
rect 722 21814 1000 21870
rect 0 21738 1000 21814
rect 0 21682 666 21738
rect 722 21682 1000 21738
rect 0 21606 1000 21682
rect 0 21550 666 21606
rect 722 21550 1000 21606
rect 0 21474 1000 21550
rect 0 21418 666 21474
rect 722 21418 1000 21474
rect 0 21342 1000 21418
rect 0 21286 666 21342
rect 722 21286 1000 21342
rect 0 21210 1000 21286
rect 0 21154 666 21210
rect 722 21154 1000 21210
rect 0 21078 1000 21154
rect 0 21022 666 21078
rect 722 21022 1000 21078
rect 0 20946 1000 21022
rect 0 20890 666 20946
rect 722 20890 1000 20946
rect 0 20814 1000 20890
rect 0 20758 666 20814
rect 722 20758 1000 20814
rect 0 20682 1000 20758
rect 0 20626 666 20682
rect 722 20626 1000 20682
rect 0 20400 1000 20626
rect 0 19978 1000 20200
rect 0 19922 666 19978
rect 722 19922 1000 19978
rect 0 19846 1000 19922
rect 0 19790 666 19846
rect 722 19790 1000 19846
rect 0 19714 1000 19790
rect 0 19658 666 19714
rect 722 19658 1000 19714
rect 0 19582 1000 19658
rect 0 19526 666 19582
rect 722 19526 1000 19582
rect 0 19450 1000 19526
rect 0 19394 666 19450
rect 722 19394 1000 19450
rect 0 19318 1000 19394
rect 0 19262 666 19318
rect 722 19262 1000 19318
rect 0 19186 1000 19262
rect 0 19130 666 19186
rect 722 19130 1000 19186
rect 0 19054 1000 19130
rect 0 18998 666 19054
rect 722 18998 1000 19054
rect 0 18922 1000 18998
rect 0 18866 666 18922
rect 722 18866 1000 18922
rect 0 18790 1000 18866
rect 0 18734 666 18790
rect 722 18734 1000 18790
rect 0 18658 1000 18734
rect 0 18602 666 18658
rect 722 18602 1000 18658
rect 0 18526 1000 18602
rect 0 18470 666 18526
rect 722 18470 1000 18526
rect 0 18394 1000 18470
rect 0 18338 666 18394
rect 722 18338 1000 18394
rect 0 18262 1000 18338
rect 0 18206 666 18262
rect 722 18206 1000 18262
rect 0 18130 1000 18206
rect 0 18074 666 18130
rect 722 18074 1000 18130
rect 0 17998 1000 18074
rect 0 17942 666 17998
rect 722 17942 1000 17998
rect 0 17866 1000 17942
rect 0 17810 666 17866
rect 722 17810 1000 17866
rect 0 17734 1000 17810
rect 0 17678 666 17734
rect 722 17678 1000 17734
rect 0 17602 1000 17678
rect 0 17546 666 17602
rect 722 17546 1000 17602
rect 0 17470 1000 17546
rect 0 17414 666 17470
rect 722 17414 1000 17470
rect 0 17200 1000 17414
rect 0 16778 1000 17000
rect 0 16722 666 16778
rect 722 16722 1000 16778
rect 0 16646 1000 16722
rect 0 16590 666 16646
rect 722 16590 1000 16646
rect 0 16514 1000 16590
rect 0 16458 666 16514
rect 722 16458 1000 16514
rect 0 16382 1000 16458
rect 0 16326 666 16382
rect 722 16326 1000 16382
rect 0 16250 1000 16326
rect 0 16194 666 16250
rect 722 16194 1000 16250
rect 0 16118 1000 16194
rect 0 16062 666 16118
rect 722 16062 1000 16118
rect 0 15986 1000 16062
rect 0 15930 666 15986
rect 722 15930 1000 15986
rect 0 15854 1000 15930
rect 0 15798 666 15854
rect 722 15798 1000 15854
rect 0 15722 1000 15798
rect 0 15666 666 15722
rect 722 15666 1000 15722
rect 0 15590 1000 15666
rect 0 15534 666 15590
rect 722 15534 1000 15590
rect 0 15458 1000 15534
rect 0 15402 666 15458
rect 722 15402 1000 15458
rect 0 15326 1000 15402
rect 0 15270 666 15326
rect 722 15270 1000 15326
rect 0 15194 1000 15270
rect 0 15138 666 15194
rect 722 15138 1000 15194
rect 0 15062 1000 15138
rect 0 15006 666 15062
rect 722 15006 1000 15062
rect 0 14930 1000 15006
rect 0 14874 666 14930
rect 722 14874 1000 14930
rect 0 14798 1000 14874
rect 0 14742 666 14798
rect 722 14742 1000 14798
rect 0 14666 1000 14742
rect 0 14610 666 14666
rect 722 14610 1000 14666
rect 0 14534 1000 14610
rect 0 14478 666 14534
rect 722 14478 1000 14534
rect 0 14402 1000 14478
rect 0 14346 666 14402
rect 722 14346 1000 14402
rect 0 14270 1000 14346
rect 0 14214 666 14270
rect 722 14214 1000 14270
rect 0 14000 1000 14214
use M1_PSUB_CDNS_40661956134174  M1_PSUB_CDNS_40661956134174_0
timestamp 1666464484
transform 1 0 500 0 -1 13192
box 0 0 1 1
use M1_PSUB_CDNS_40661956134174  M1_PSUB_CDNS_40661956134174_1
timestamp 1666464484
transform 1 0 500 0 1 69873
box 0 0 1 1
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_0
timestamp 1666464484
transform -1 0 48 0 1 41524
box 0 0 1 1
use M1_PSUB_CDNS_40661956134176  M1_PSUB_CDNS_40661956134176_1
timestamp 1666464484
transform 1 0 952 0 1 41524
box 0 0 1 1
use M2_M1_CDNS_40661956134173  M2_M1_CDNS_40661956134173_0
timestamp 1666464484
transform 1 0 877 0 1 49900
box 0 0 1 1
use M2_M1_CDNS_40661956134173  M2_M1_CDNS_40661956134173_1
timestamp 1666464484
transform 1 0 877 0 1 64300
box 0 0 1 1
use M2_M1_CDNS_40661956134173  M2_M1_CDNS_40661956134173_2
timestamp 1666464484
transform 1 0 85 0 1 64300
box 0 0 1 1
use M2_M1_CDNS_40661956134173  M2_M1_CDNS_40661956134173_3
timestamp 1666464484
transform 1 0 85 0 1 49900
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_0
timestamp 1666464484
transform 1 0 510 0 1 62697
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_1
timestamp 1666464484
transform 1 0 694 0 1 69023
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_2
timestamp 1666464484
transform 1 0 694 0 1 65910
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_3
timestamp 1666464484
transform 1 0 318 0 1 67494
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_4
timestamp 1666464484
transform 1 0 694 0 1 61108
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_5
timestamp 1666464484
transform 1 0 694 0 1 57897
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_6
timestamp 1666464484
transform 1 0 694 0 1 40327
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_7
timestamp 1666464484
transform 1 0 318 0 1 59505
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_8
timestamp 1666464484
transform 1 0 318 0 1 56323
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_9
timestamp 1666464484
transform 1 0 318 0 1 54704
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_10
timestamp 1666464484
transform 1 0 318 0 1 53113
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_11
timestamp 1666464484
transform 1 0 318 0 1 41895
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_12
timestamp 1666464484
transform 1 0 318 0 1 24298
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_13
timestamp 1666464484
transform 1 0 510 0 1 51504
box 0 0 1 1
use M3_M2_CDNS_40661956134172  M3_M2_CDNS_40661956134172_14
timestamp 1666464484
transform 1 0 694 0 1 25929
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_0
timestamp 1666464484
transform 1 0 694 0 1 47528
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_1
timestamp 1666464484
transform 1 0 694 0 1 21908
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_2
timestamp 1666464484
transform 1 0 694 0 1 15496
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_3
timestamp 1666464484
transform 1 0 318 0 1 44311
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_4
timestamp 1666464484
transform 1 0 318 0 1 37888
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_5
timestamp 1666464484
transform 1 0 318 0 1 34718
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_6
timestamp 1666464484
transform 1 0 318 0 1 31513
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_7
timestamp 1666464484
transform 1 0 318 0 1 28343
box 0 0 1 1
use M3_M2_CDNS_40661956134175  M3_M2_CDNS_40661956134175_8
timestamp 1666464484
transform 1 0 694 0 1 18696
box 0 0 1 1
use M3_M2_CDNS_40661956134177  M3_M2_CDNS_40661956134177_0
timestamp 1666464484
transform 1 0 85 0 1 49900
box 0 0 1 1
use M3_M2_CDNS_40661956134177  M3_M2_CDNS_40661956134177_1
timestamp 1666464484
transform 1 0 877 0 1 64300
box 0 0 1 1
use M3_M2_CDNS_40661956134177  M3_M2_CDNS_40661956134177_2
timestamp 1666464484
transform 1 0 85 0 1 64300
box 0 0 1 1
use M3_M2_CDNS_40661956134177  M3_M2_CDNS_40661956134177_3
timestamp 1666464484
transform 1 0 877 0 1 49900
box 0 0 1 1
use POLY_SUB_FILL  POLY_SUB_FILL_0
array 0 0 0 0 34 1600
timestamp 1666464484
transform 1 0 -806 0 1 13819
box 880 -349 1727 1343
<< labels >>
rlabel metal3 s 800 49200 1000 50600 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 63600 1000 65000 4 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 800 50800 1000 52200 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 62000 1000 63400 4 VDD
port 3 nsew power bidirectional
rlabel metal3 s 800 14000 1000 17000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 17200 1000 20200 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 20400 1000 23400 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 46000 1000 49000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 25200 1000 26600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 39600 1000 41000 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 57200 1000 58600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 60400 1000 61800 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 65200 1000 66600 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 68400 1000 69678 4 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 800 26800 1000 29800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 30000 1000 33000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 33200 1000 36200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 36400 1000 39400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 42800 1000 45800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 23600 1000 25000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 41200 1000 42600 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 52400 1000 53800 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 54000 1000 55400 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 55600 1000 57000 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 58800 1000 60200 4 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 800 66800 1000 68200 4 DVDD
port 1 nsew power bidirectional
rlabel space 0 400 0 400 4 & Metric 1.00
rlabel space 0 800 0 800 4 & Version 2014q3v1
rlabel space 0 1200 0 1200 4 & Product GF018green_ipio_5p0c_75
rlabel space 0 1600 0 1600 4 & Vendor GLOBALFOUNDRIES
rlabel metal3 s 0 66800 200 68200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 58800 200 60200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 55600 200 57000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 54000 200 55400 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 52400 200 53800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 42800 200 45800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 41200 200 42600 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 36400 200 39400 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 33200 200 36200 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 30000 200 33000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 26800 200 29800 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 23600 200 25000 1 DVDD
port 1 nsew power bidirectional
rlabel metal3 s 0 68400 200 69678 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 65200 200 66600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 60400 200 61800 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 57200 200 58600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 46000 200 49000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 39600 200 41000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 25200 200 26600 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 20400 200 23400 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 17200 200 20200 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 14000 200 17000 1 DVSS
port 2 nsew ground bidirectional
rlabel metal3 s 0 62000 200 63400 1 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 50800 200 52200 1 VDD
port 3 nsew power bidirectional
rlabel metal3 s 0 63600 200 65000 1 VSS
port 4 nsew ground bidirectional
rlabel metal3 s 0 49200 200 50600 1 VSS
port 4 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 1000 70000
string GDS_END 4162130
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 4155950
string LEFclass PAD SPACER
string LEFsite GF_IO_Site
string LEFsymmetry X Y R90
<< end >>
