magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 352 4118 870
<< pwell >>
rect -86 -86 4118 352
<< mvnmos >>
rect 179 68 299 140
rect 403 68 523 140
rect 571 68 691 140
rect 1027 68 1147 140
rect 1195 68 1315 140
rect 1419 68 1539 140
rect 1587 68 1707 140
rect 2083 68 2203 140
rect 2251 68 2371 140
rect 2475 68 2595 140
rect 2643 68 2763 140
rect 3119 68 3239 141
rect 3287 68 3407 141
rect 3547 68 3667 232
rect 3771 68 3891 232
<< mvpmos >>
rect 179 644 279 716
rect 403 644 503 716
rect 571 644 671 716
rect 1007 644 1107 716
rect 1175 644 1275 716
rect 1459 644 1559 716
rect 1627 644 1727 716
rect 2063 644 2163 716
rect 2231 644 2331 716
rect 2515 644 2615 716
rect 2683 644 2783 716
rect 3119 622 3219 694
rect 3287 622 3387 694
rect 3567 472 3667 716
rect 3771 472 3871 716
<< mvndiff >>
rect 47 180 119 193
rect 47 134 60 180
rect 106 140 119 180
rect 751 200 823 213
rect 751 154 764 200
rect 810 154 823 200
rect 751 140 823 154
rect 106 134 179 140
rect 47 68 179 134
rect 299 127 403 140
rect 299 81 328 127
rect 374 81 403 127
rect 299 68 403 81
rect 523 68 571 140
rect 691 68 823 140
rect 895 200 967 213
rect 895 154 908 200
rect 954 154 967 200
rect 895 140 967 154
rect 1767 200 1839 213
rect 1767 154 1780 200
rect 1826 154 1839 200
rect 1767 140 1839 154
rect 895 68 1027 140
rect 1147 68 1195 140
rect 1315 127 1419 140
rect 1315 81 1344 127
rect 1390 81 1419 127
rect 1315 68 1419 81
rect 1539 68 1587 140
rect 1707 68 1839 140
rect 1951 200 2023 213
rect 1951 154 1964 200
rect 2010 154 2023 200
rect 1951 140 2023 154
rect 2823 200 2895 213
rect 2823 154 2836 200
rect 2882 154 2895 200
rect 2823 140 2895 154
rect 1951 68 2083 140
rect 2203 68 2251 140
rect 2371 127 2475 140
rect 2371 81 2400 127
rect 2446 81 2475 127
rect 2371 68 2475 81
rect 2595 68 2643 140
rect 2763 68 2895 140
rect 2987 200 3059 213
rect 2987 154 3000 200
rect 3046 154 3059 200
rect 2987 141 3059 154
rect 3467 141 3547 232
rect 2987 68 3119 141
rect 3239 68 3287 141
rect 3407 127 3547 141
rect 3407 81 3436 127
rect 3482 81 3547 127
rect 3407 68 3547 81
rect 3667 192 3771 232
rect 3667 146 3696 192
rect 3742 146 3771 192
rect 3667 68 3771 146
rect 3891 127 3979 232
rect 3891 81 3920 127
rect 3966 81 3979 127
rect 3891 68 3979 81
<< mvpdiff >>
rect 47 644 179 716
rect 279 703 403 716
rect 279 657 308 703
rect 354 657 403 703
rect 279 644 403 657
rect 503 644 571 716
rect 671 644 803 716
rect 47 621 119 644
rect 47 575 60 621
rect 106 575 119 621
rect 47 562 119 575
rect 731 621 803 644
rect 731 575 744 621
rect 790 575 803 621
rect 731 562 803 575
rect 875 644 1007 716
rect 1107 644 1175 716
rect 1275 703 1459 716
rect 1275 657 1304 703
rect 1350 657 1459 703
rect 1275 644 1459 657
rect 1559 644 1627 716
rect 1727 644 1859 716
rect 875 621 947 644
rect 875 575 888 621
rect 934 575 947 621
rect 875 562 947 575
rect 1787 621 1859 644
rect 1787 575 1800 621
rect 1846 575 1859 621
rect 1787 562 1859 575
rect 1931 644 2063 716
rect 2163 644 2231 716
rect 2331 703 2515 716
rect 2331 657 2360 703
rect 2406 657 2515 703
rect 2331 644 2515 657
rect 2615 644 2683 716
rect 2783 644 2915 716
rect 3447 694 3567 716
rect 1931 621 2003 644
rect 1931 575 1944 621
rect 1990 575 2003 621
rect 1931 562 2003 575
rect 2843 621 2915 644
rect 2843 575 2856 621
rect 2902 575 2915 621
rect 2843 562 2915 575
rect 2987 622 3119 694
rect 3219 622 3287 694
rect 3387 665 3567 694
rect 3387 622 3492 665
rect 2987 621 3059 622
rect 2987 575 3000 621
rect 3046 575 3059 621
rect 2987 562 3059 575
rect 3447 525 3492 622
rect 3538 525 3567 665
rect 3447 472 3567 525
rect 3667 665 3771 716
rect 3667 525 3696 665
rect 3742 525 3771 665
rect 3667 472 3771 525
rect 3871 665 3959 716
rect 3871 525 3900 665
rect 3946 525 3959 665
rect 3871 472 3959 525
<< mvndiffc >>
rect 60 134 106 180
rect 764 154 810 200
rect 328 81 374 127
rect 908 154 954 200
rect 1780 154 1826 200
rect 1344 81 1390 127
rect 1964 154 2010 200
rect 2836 154 2882 200
rect 2400 81 2446 127
rect 3000 154 3046 200
rect 3436 81 3482 127
rect 3696 146 3742 192
rect 3920 81 3966 127
<< mvpdiffc >>
rect 308 657 354 703
rect 60 575 106 621
rect 744 575 790 621
rect 1304 657 1350 703
rect 888 575 934 621
rect 1800 575 1846 621
rect 2360 657 2406 703
rect 1944 575 1990 621
rect 2856 575 2902 621
rect 3000 575 3046 621
rect 3492 525 3538 665
rect 3696 525 3742 665
rect 3900 525 3946 665
<< polysilicon >>
rect 179 716 279 760
rect 403 716 503 760
rect 571 716 671 760
rect 1007 716 1107 760
rect 1175 716 1275 760
rect 1459 716 1559 760
rect 1627 716 1727 760
rect 2063 716 2163 760
rect 2231 716 2331 760
rect 2515 716 2615 760
rect 2683 716 2783 760
rect 179 303 279 644
rect 179 257 192 303
rect 238 257 279 303
rect 179 184 279 257
rect 403 483 503 644
rect 571 483 671 644
rect 403 470 671 483
rect 403 424 416 470
rect 462 424 596 470
rect 642 424 671 470
rect 403 411 671 424
rect 403 184 503 411
rect 571 184 671 411
rect 1007 371 1107 644
rect 1175 371 1275 644
rect 1007 350 1275 371
rect 1007 304 1020 350
rect 1066 304 1275 350
rect 1007 290 1275 304
rect 179 140 299 184
rect 403 140 523 184
rect 571 140 691 184
rect 1027 140 1147 290
rect 1195 184 1275 290
rect 1459 371 1559 644
rect 1627 371 1727 644
rect 3119 694 3219 738
rect 3287 694 3387 738
rect 3567 716 3667 760
rect 3771 716 3871 760
rect 1459 350 1727 371
rect 1459 304 1472 350
rect 1612 304 1727 350
rect 1459 290 1727 304
rect 2063 371 2163 644
rect 2231 371 2331 644
rect 2063 350 2331 371
rect 2063 304 2076 350
rect 2122 304 2331 350
rect 2063 290 2331 304
rect 1459 184 1539 290
rect 1195 140 1315 184
rect 1419 140 1539 184
rect 1587 140 1707 290
rect 2083 140 2203 290
rect 2251 184 2331 290
rect 2515 371 2615 644
rect 2683 371 2783 644
rect 2515 350 2783 371
rect 2515 304 2528 350
rect 2668 304 2783 350
rect 2515 290 2783 304
rect 3119 377 3219 622
rect 3287 377 3387 622
rect 3119 364 3387 377
rect 3119 318 3132 364
rect 3272 318 3387 364
rect 3567 340 3667 472
rect 3771 340 3871 472
rect 3567 325 3891 340
rect 3567 323 3580 325
rect 3119 305 3387 318
rect 2515 184 2595 290
rect 2251 140 2371 184
rect 2475 140 2595 184
rect 2643 140 2763 290
rect 3119 185 3219 305
rect 3287 185 3387 305
rect 3547 279 3580 323
rect 3626 292 3891 325
rect 3626 279 3667 292
rect 3547 232 3667 279
rect 3771 232 3891 292
rect 3119 141 3239 185
rect 3287 141 3407 185
rect 179 24 299 68
rect 403 24 523 68
rect 571 24 691 68
rect 1027 24 1147 68
rect 1195 24 1315 68
rect 1419 24 1539 68
rect 1587 24 1707 68
rect 2083 24 2203 68
rect 2251 24 2371 68
rect 2475 24 2595 68
rect 2643 24 2763 68
rect 3119 24 3239 68
rect 3287 24 3407 68
rect 3547 24 3667 68
rect 3771 24 3891 68
<< polycontact >>
rect 192 257 238 303
rect 416 424 462 470
rect 596 424 642 470
rect 1020 304 1066 350
rect 1472 304 1612 350
rect 2076 304 2122 350
rect 2528 304 2668 350
rect 3132 318 3272 364
rect 3580 279 3626 325
<< metal1 >>
rect 0 724 4032 844
rect 297 703 365 724
rect 297 657 308 703
rect 354 657 365 703
rect 1293 703 1361 724
rect 1293 657 1304 703
rect 1350 657 1361 703
rect 2349 703 2417 724
rect 2349 657 2360 703
rect 2406 657 2417 703
rect 3492 665 3538 724
rect 744 621 790 632
rect 1780 621 1857 632
rect 2836 621 2913 632
rect 49 575 60 621
rect 106 575 117 621
rect 49 481 117 575
rect 877 575 888 621
rect 934 575 1158 621
rect 49 470 653 481
rect 49 424 416 470
rect 462 424 596 470
rect 642 424 653 470
rect 49 413 653 424
rect 49 180 95 413
rect 744 361 790 575
rect 744 350 1066 361
rect 186 303 679 320
rect 186 257 192 303
rect 238 257 679 303
rect 186 240 679 257
rect 744 304 1020 350
rect 744 293 1066 304
rect 1112 350 1158 575
rect 1780 575 1800 621
rect 1846 575 1857 621
rect 1933 575 1944 621
rect 1990 575 2214 621
rect 1780 564 1857 575
rect 1780 361 1826 564
rect 1780 350 2122 361
rect 1112 304 1472 350
rect 1612 304 1623 350
rect 1780 304 2076 350
rect 744 200 821 293
rect 1112 200 1158 304
rect 49 134 60 180
rect 106 134 117 180
rect 744 154 764 200
rect 810 154 821 200
rect 897 154 908 200
rect 954 154 1158 200
rect 1780 293 2122 304
rect 2168 350 2214 575
rect 2836 575 2856 621
rect 2902 575 2913 621
rect 2836 564 2913 575
rect 3000 621 3046 632
rect 2836 375 2882 564
rect 3000 493 3046 575
rect 3492 506 3538 525
rect 3696 665 3790 676
rect 3742 525 3790 665
rect 3000 447 3376 493
rect 2836 364 3272 375
rect 2168 304 2528 350
rect 2668 304 2679 350
rect 2836 318 3132 364
rect 2836 307 3272 318
rect 3330 325 3376 447
rect 1780 200 1826 293
rect 2168 200 2214 304
rect 1953 154 1964 200
rect 2010 154 2214 200
rect 2836 200 2882 307
rect 3330 279 3580 325
rect 3626 279 3637 325
rect 3330 200 3376 279
rect 2989 154 3000 200
rect 3046 154 3376 200
rect 3696 192 3790 525
rect 3900 665 3946 724
rect 3900 506 3946 525
rect 1780 143 1826 154
rect 2836 143 2882 154
rect 3742 146 3790 192
rect 3436 127 3482 138
rect 3696 135 3790 146
rect 317 81 328 127
rect 374 81 385 127
rect 317 60 385 81
rect 1333 81 1344 127
rect 1390 81 1401 127
rect 1333 60 1401 81
rect 2389 81 2400 127
rect 2446 81 2457 127
rect 2389 60 2457 81
rect 3436 60 3482 81
rect 3920 127 3966 138
rect 3920 60 3966 81
rect 0 -60 4032 60
<< labels >>
flabel metal1 s 0 724 4032 844 0 FreeSans 400 0 0 0 VDD
port 3 nsew power bidirectional abutment
flabel metal1 s 186 240 679 320 0 FreeSans 400 0 0 0 I
port 1 nsew default input
flabel metal1 s 3920 127 3966 138 0 FreeSans 400 0 0 0 VSS
port 6 nsew ground bidirectional abutment
flabel metal1 s 3696 135 3790 676 0 FreeSans 400 0 0 0 Z
port 2 nsew default output
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 3900 657 3946 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3492 657 3538 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 2349 657 2417 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 1293 657 1361 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 297 657 365 724 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3900 506 3946 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3492 506 3538 657 1 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 3436 127 3482 138 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3920 60 3966 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 3436 60 3482 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 2389 60 2457 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 1333 60 1401 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 317 60 385 127 1 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4032 60 1 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4032 784
string GDS_END 1114712
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1107668
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
