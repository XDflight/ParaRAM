magic
tech gf180mcuA
timestamp 1666464484
<< properties >>
string GDS_END 518674
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 493966
<< end >>
