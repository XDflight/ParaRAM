magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -144 -4186 1106 -3712
<< nmos >>
rect 197 -10182 317 -7687
rect 421 -10182 541 -7687
rect 645 -10182 765 -7687
<< ndiff >>
rect 78 -7733 197 -7687
rect 78 -7779 122 -7733
rect 168 -7779 197 -7733
rect 78 -7900 197 -7779
rect 78 -7946 122 -7900
rect 168 -7946 197 -7900
rect 78 -8068 197 -7946
rect 78 -8114 122 -8068
rect 168 -8114 197 -8068
rect 78 -8236 197 -8114
rect 78 -8282 122 -8236
rect 168 -8282 197 -8236
rect 78 -8404 197 -8282
rect 78 -8450 122 -8404
rect 168 -8450 197 -8404
rect 78 -8571 197 -8450
rect 78 -8617 122 -8571
rect 168 -8617 197 -8571
rect 78 -8739 197 -8617
rect 78 -8785 122 -8739
rect 168 -8785 197 -8739
rect 78 -8907 197 -8785
rect 78 -8953 122 -8907
rect 168 -8953 197 -8907
rect 78 -9075 197 -8953
rect 78 -9121 122 -9075
rect 168 -9121 197 -9075
rect 78 -9243 197 -9121
rect 78 -9289 122 -9243
rect 168 -9289 197 -9243
rect 78 -9410 197 -9289
rect 78 -9456 122 -9410
rect 168 -9456 197 -9410
rect 78 -9580 197 -9456
rect 78 -9626 122 -9580
rect 168 -9626 197 -9580
rect 78 -9750 197 -9626
rect 78 -9796 122 -9750
rect 168 -9796 197 -9750
rect 78 -9920 197 -9796
rect 78 -9966 122 -9920
rect 168 -9966 197 -9920
rect 78 -10090 197 -9966
rect 78 -10136 122 -10090
rect 168 -10136 197 -10090
rect 78 -10182 197 -10136
rect 317 -10182 421 -7687
rect 541 -10182 645 -7687
rect 765 -7733 883 -7687
rect 765 -7779 794 -7733
rect 840 -7779 883 -7733
rect 765 -7900 883 -7779
rect 765 -7946 794 -7900
rect 840 -7946 883 -7900
rect 765 -8068 883 -7946
rect 765 -8114 794 -8068
rect 840 -8114 883 -8068
rect 765 -8236 883 -8114
rect 765 -8282 794 -8236
rect 840 -8282 883 -8236
rect 765 -8404 883 -8282
rect 765 -8450 794 -8404
rect 840 -8450 883 -8404
rect 765 -8571 883 -8450
rect 765 -8617 794 -8571
rect 840 -8617 883 -8571
rect 765 -8739 883 -8617
rect 765 -8785 794 -8739
rect 840 -8785 883 -8739
rect 765 -8907 883 -8785
rect 765 -8953 794 -8907
rect 840 -8953 883 -8907
rect 765 -9075 883 -8953
rect 765 -9121 794 -9075
rect 840 -9121 883 -9075
rect 765 -9243 883 -9121
rect 765 -9289 794 -9243
rect 840 -9289 883 -9243
rect 765 -9410 883 -9289
rect 765 -9456 794 -9410
rect 840 -9456 883 -9410
rect 765 -9580 883 -9456
rect 765 -9626 794 -9580
rect 840 -9626 883 -9580
rect 765 -9750 883 -9626
rect 765 -9796 794 -9750
rect 840 -9796 883 -9750
rect 765 -9920 883 -9796
rect 765 -9966 794 -9920
rect 840 -9966 883 -9920
rect 765 -10090 883 -9966
rect 765 -10136 794 -10090
rect 840 -10136 883 -10090
rect 765 -10182 883 -10136
<< ndiffc >>
rect 122 -7779 168 -7733
rect 122 -7946 168 -7900
rect 122 -8114 168 -8068
rect 122 -8282 168 -8236
rect 122 -8450 168 -8404
rect 122 -8617 168 -8571
rect 122 -8785 168 -8739
rect 122 -8953 168 -8907
rect 122 -9121 168 -9075
rect 122 -9289 168 -9243
rect 122 -9456 168 -9410
rect 122 -9626 168 -9580
rect 122 -9796 168 -9750
rect 122 -9966 168 -9920
rect 122 -10136 168 -10090
rect 794 -7779 840 -7733
rect 794 -7946 840 -7900
rect 794 -8114 840 -8068
rect 794 -8282 840 -8236
rect 794 -8450 840 -8404
rect 794 -8617 840 -8571
rect 794 -8785 840 -8739
rect 794 -8953 840 -8907
rect 794 -9121 840 -9075
rect 794 -9289 840 -9243
rect 794 -9456 840 -9410
rect 794 -9626 840 -9580
rect 794 -9796 840 -9750
rect 794 -9966 840 -9920
rect 794 -10136 840 -10090
<< psubdiff >>
rect -1 186 963 245
rect -1 140 212 186
rect 258 140 370 186
rect 416 140 528 186
rect 574 140 686 186
rect 732 140 963 186
rect -1 81 963 140
rect -1 -10458 963 -10399
rect -1 -10504 212 -10458
rect 258 -10504 370 -10458
rect 416 -10504 528 -10458
rect 574 -10504 686 -10458
rect 732 -10504 963 -10458
rect -1 -10563 963 -10504
<< nsubdiff >>
rect -1 -3935 963 -3879
rect -1 -3981 201 -3935
rect 247 -3981 359 -3935
rect 405 -3981 517 -3935
rect 563 -3981 963 -3935
rect -1 -4039 963 -3981
<< psubdiffcont >>
rect 212 140 258 186
rect 370 140 416 186
rect 528 140 574 186
rect 686 140 732 186
rect 212 -10504 258 -10458
rect 370 -10504 416 -10458
rect 528 -10504 574 -10458
rect 686 -10504 732 -10458
<< nsubdiffcont >>
rect 201 -3981 247 -3935
rect 359 -3981 405 -3935
rect 517 -3981 563 -3935
<< polysilicon >>
rect 197 -1115 317 -1074
rect 421 -1115 541 -1074
rect 645 -1115 765 -1074
rect 197 -1252 765 -1115
rect 197 -1311 317 -1252
rect 421 -1311 541 -1252
rect 645 -1311 765 -1252
rect 197 -3654 317 -3627
rect 421 -3654 541 -3634
rect 645 -3654 765 -3634
rect 197 -3698 765 -3654
rect 197 -3744 327 -3698
rect 655 -3744 765 -3698
rect 197 -3791 765 -3744
rect 197 -6820 317 -6353
rect 197 -6957 318 -6820
rect 197 -7687 317 -6957
rect 421 -7687 541 -6353
rect 645 -7687 765 -6353
rect 197 -10255 317 -10182
rect 421 -10255 541 -10182
rect 645 -10255 765 -10182
<< polycontact >>
rect 327 -3744 655 -3698
<< metal1 >>
rect -1 186 963 236
rect -1 140 212 186
rect 258 140 370 186
rect 416 140 528 186
rect 574 167 686 186
rect -1 115 574 140
rect 626 140 686 167
rect 732 140 963 186
rect 626 115 963 140
rect -1 -51 963 115
rect -1 -55 574 -51
rect 87 -56 203 -55
rect 87 -250 202 -56
rect 535 -103 574 -55
rect 626 -55 963 -51
rect 626 -103 664 -55
rect 303 -184 431 -145
rect 303 -236 341 -184
rect 393 -236 431 -184
rect 303 -402 431 -236
rect 535 -250 664 -103
rect 303 -454 341 -402
rect 393 -454 431 -402
rect 303 -620 431 -454
rect 536 -269 664 -250
rect 536 -321 574 -269
rect 626 -321 664 -269
rect 536 -487 664 -321
rect 536 -539 574 -487
rect 626 -539 664 -487
rect 536 -579 664 -539
rect 303 -672 341 -620
rect 393 -672 431 -620
rect 303 -712 431 -672
rect 311 -1120 426 -960
rect 759 -1120 874 -960
rect 311 -1239 874 -1120
rect 311 -1240 427 -1239
rect 311 -1384 426 -1240
rect 759 -1384 874 -1239
rect 81 -2925 209 -2886
rect 81 -2977 119 -2925
rect 171 -2977 209 -2925
rect 81 -3143 209 -2977
rect 81 -3195 119 -3143
rect 171 -3195 209 -3143
rect 81 -3361 209 -3195
rect 81 -3413 119 -3361
rect 171 -3413 209 -3361
rect 81 -3453 209 -3413
rect 529 -2925 657 -2886
rect 529 -2977 567 -2925
rect 619 -2977 657 -2925
rect 529 -3143 657 -2977
rect 529 -3195 567 -3143
rect 619 -3195 657 -3143
rect 529 -3361 657 -3195
rect 529 -3413 567 -3361
rect 619 -3413 657 -3361
rect 529 -3453 657 -3413
rect 199 -3698 874 -3663
rect 199 -3744 327 -3698
rect 655 -3744 874 -3698
rect 199 -3782 874 -3744
rect -1 -3935 650 -3899
rect -1 -3981 201 -3935
rect 247 -3981 359 -3935
rect 405 -3981 517 -3935
rect 563 -3981 650 -3935
rect -1 -4006 650 -3981
rect -1 -4018 653 -4006
rect 81 -4045 209 -4018
rect 81 -4097 119 -4045
rect 171 -4097 209 -4045
rect 81 -4263 209 -4097
rect 81 -4315 119 -4263
rect 171 -4315 209 -4263
rect 81 -4480 209 -4315
rect 81 -4532 119 -4480
rect 171 -4532 209 -4480
rect 81 -4698 209 -4532
rect 81 -4750 119 -4698
rect 171 -4750 209 -4698
rect 81 -4916 209 -4750
rect 81 -4968 119 -4916
rect 171 -4968 209 -4916
rect 81 -5133 209 -4968
rect 81 -5185 119 -5133
rect 171 -5185 209 -5133
rect 81 -5351 209 -5185
rect 81 -5403 119 -5351
rect 171 -5403 209 -5351
rect 81 -5443 209 -5403
rect 525 -4045 653 -4018
rect 525 -4097 563 -4045
rect 615 -4097 653 -4045
rect 525 -4263 653 -4097
rect 525 -4315 563 -4263
rect 615 -4315 653 -4263
rect 525 -4480 653 -4315
rect 759 -4333 874 -3782
rect 525 -4532 563 -4480
rect 615 -4532 653 -4480
rect 525 -4698 653 -4532
rect 525 -4750 563 -4698
rect 615 -4750 653 -4698
rect 525 -4916 653 -4750
rect 525 -4968 563 -4916
rect 615 -4968 653 -4916
rect 525 -5133 653 -4968
rect 525 -5185 563 -5133
rect 615 -5185 653 -5133
rect 525 -5351 653 -5185
rect 525 -5403 563 -5351
rect 615 -5403 653 -5351
rect 525 -5443 653 -5403
rect 94 -5444 209 -5443
rect 538 -5444 653 -5443
rect 307 -5995 431 -5955
rect 307 -6047 343 -5995
rect 395 -6047 431 -5995
rect 307 -6213 431 -6047
rect 307 -6265 343 -6213
rect 395 -6265 431 -6213
rect 307 -6305 431 -6265
rect 755 -5995 879 -5955
rect 755 -6047 791 -5995
rect 843 -6047 879 -5995
rect 755 -6213 879 -6047
rect 755 -6265 791 -6213
rect 843 -6265 879 -6213
rect 755 -6305 879 -6265
rect -58 -6530 1020 -6438
rect -58 -6732 1020 -6640
rect -58 -6933 1020 -6842
rect -58 -7135 1020 -7043
rect -58 -7337 1020 -7245
rect -58 -7539 1020 -7447
rect 87 -7733 202 -7696
rect 87 -7779 122 -7733
rect 168 -7779 202 -7733
rect 87 -7801 202 -7779
rect 759 -7733 875 -7696
rect 759 -7779 794 -7733
rect 840 -7779 875 -7733
rect 87 -7900 203 -7801
rect 87 -7946 122 -7900
rect 168 -7946 203 -7900
rect 87 -8068 203 -7946
rect 87 -8114 122 -8068
rect 168 -8114 203 -8068
rect 87 -8236 203 -8114
rect 87 -8282 122 -8236
rect 168 -8282 203 -8236
rect 87 -8404 203 -8282
rect 87 -8450 122 -8404
rect 168 -8450 203 -8404
rect 87 -8571 203 -8450
rect 87 -8617 122 -8571
rect 168 -8617 203 -8571
rect 87 -8739 203 -8617
rect 87 -8785 122 -8739
rect 168 -8785 203 -8739
rect 87 -8907 203 -8785
rect 87 -8953 122 -8907
rect 168 -8953 203 -8907
rect 87 -9075 203 -8953
rect 87 -9121 122 -9075
rect 168 -9121 203 -9075
rect 87 -9243 203 -9121
rect 87 -9289 122 -9243
rect 168 -9289 203 -9243
rect 87 -9410 203 -9289
rect 87 -9456 122 -9410
rect 168 -9456 203 -9410
rect 87 -9580 203 -9456
rect 87 -9626 122 -9580
rect 168 -9626 203 -9580
rect 87 -9750 203 -9626
rect 87 -9796 122 -9750
rect 168 -9796 203 -9750
rect 87 -9920 203 -9796
rect 87 -9966 122 -9920
rect 168 -9966 203 -9920
rect 87 -10090 203 -9966
rect 87 -10136 122 -10090
rect 168 -10136 203 -10090
rect 87 -10262 203 -10136
rect 759 -7900 875 -7779
rect 759 -7946 794 -7900
rect 840 -7946 875 -7900
rect 759 -8068 875 -7946
rect 759 -8114 794 -8068
rect 840 -8114 875 -8068
rect 759 -8236 875 -8114
rect 759 -8282 794 -8236
rect 840 -8282 875 -8236
rect 759 -8404 875 -8282
rect 759 -8450 794 -8404
rect 840 -8450 875 -8404
rect 759 -8571 875 -8450
rect 759 -8617 794 -8571
rect 840 -8617 875 -8571
rect 759 -8739 875 -8617
rect 759 -8785 794 -8739
rect 840 -8785 875 -8739
rect 759 -8907 875 -8785
rect 759 -8953 794 -8907
rect 840 -8953 875 -8907
rect 759 -9075 875 -8953
rect 759 -9121 794 -9075
rect 840 -9121 875 -9075
rect 759 -9243 875 -9121
rect 759 -9289 794 -9243
rect 840 -9289 875 -9243
rect 759 -9353 875 -9289
rect 759 -9410 874 -9353
rect 759 -9456 794 -9410
rect 840 -9456 874 -9410
rect 759 -9580 874 -9456
rect 759 -9626 794 -9580
rect 840 -9626 874 -9580
rect 759 -9750 874 -9626
rect 759 -9796 794 -9750
rect 840 -9796 874 -9750
rect 759 -9920 874 -9796
rect 759 -9966 794 -9920
rect 840 -9966 874 -9920
rect 759 -10090 874 -9966
rect 759 -10136 794 -10090
rect 840 -10136 874 -10090
rect 759 -10173 874 -10136
rect 81 -10263 209 -10262
rect 8 -10458 963 -10263
rect 8 -10504 212 -10458
rect 258 -10504 370 -10458
rect 416 -10504 528 -10458
rect 574 -10504 686 -10458
rect 732 -10504 963 -10458
rect 8 -10554 963 -10504
<< via1 >>
rect 574 115 626 167
rect 574 -103 626 -51
rect 341 -236 393 -184
rect 341 -454 393 -402
rect 574 -321 626 -269
rect 574 -539 626 -487
rect 341 -672 393 -620
rect 119 -2977 171 -2925
rect 119 -3195 171 -3143
rect 119 -3413 171 -3361
rect 567 -2977 619 -2925
rect 567 -3195 619 -3143
rect 567 -3413 619 -3361
rect 119 -4097 171 -4045
rect 119 -4315 171 -4263
rect 119 -4532 171 -4480
rect 119 -4750 171 -4698
rect 119 -4968 171 -4916
rect 119 -5185 171 -5133
rect 119 -5403 171 -5351
rect 563 -4097 615 -4045
rect 563 -4315 615 -4263
rect 563 -4532 615 -4480
rect 563 -4750 615 -4698
rect 563 -4968 615 -4916
rect 563 -5185 615 -5133
rect 563 -5403 615 -5351
rect 343 -6047 395 -5995
rect 343 -6265 395 -6213
rect 791 -6047 843 -5995
rect 791 -6265 843 -6213
<< metal2 >>
rect 210 -184 431 327
rect 210 -236 341 -184
rect 393 -236 431 -184
rect 210 -402 431 -236
rect 210 -454 341 -402
rect 393 -454 431 -402
rect 210 -620 431 -454
rect 536 169 664 206
rect 536 113 572 169
rect 628 113 664 169
rect 536 -49 664 113
rect 536 -105 572 -49
rect 628 -105 664 -49
rect 536 -267 664 -105
rect 536 -323 572 -267
rect 628 -323 664 -267
rect 536 -485 664 -323
rect 536 -541 572 -485
rect 628 -541 664 -485
rect 536 -579 664 -541
rect 210 -672 341 -620
rect 393 -672 431 -620
rect 210 -713 431 -672
rect 81 -2923 209 -2886
rect 81 -2979 117 -2923
rect 173 -2979 209 -2923
rect 81 -3141 209 -2979
rect 81 -3197 117 -3141
rect 173 -3197 209 -3141
rect 81 -3359 209 -3197
rect 81 -3415 117 -3359
rect 173 -3415 209 -3359
rect 81 -3453 209 -3415
rect 529 -2923 657 -2886
rect 529 -2979 565 -2923
rect 621 -2979 657 -2923
rect 529 -3141 657 -2979
rect 529 -3197 565 -3141
rect 621 -3197 657 -3141
rect 529 -3359 657 -3197
rect 529 -3415 565 -3359
rect 621 -3415 657 -3359
rect 529 -3453 657 -3415
rect 81 -4043 209 -4006
rect 81 -4099 117 -4043
rect 173 -4099 209 -4043
rect 81 -4261 209 -4099
rect 81 -4317 117 -4261
rect 173 -4317 209 -4261
rect 81 -4478 209 -4317
rect 81 -4534 117 -4478
rect 173 -4534 209 -4478
rect 81 -4696 209 -4534
rect 81 -4752 117 -4696
rect 173 -4752 209 -4696
rect 81 -4914 209 -4752
rect 81 -4970 117 -4914
rect 173 -4970 209 -4914
rect 81 -5131 209 -4970
rect 81 -5187 117 -5131
rect 173 -5187 209 -5131
rect 81 -5349 209 -5187
rect 81 -5405 117 -5349
rect 173 -5405 209 -5349
rect 81 -5443 209 -5405
rect 525 -4043 653 -4006
rect 525 -4099 561 -4043
rect 617 -4099 653 -4043
rect 525 -4261 653 -4099
rect 525 -4317 561 -4261
rect 617 -4317 653 -4261
rect 525 -4478 653 -4317
rect 525 -4534 561 -4478
rect 617 -4534 653 -4478
rect 525 -4696 653 -4534
rect 525 -4752 561 -4696
rect 617 -4752 653 -4696
rect 525 -4914 653 -4752
rect 525 -4970 561 -4914
rect 617 -4970 653 -4914
rect 525 -5131 653 -4970
rect 525 -5187 561 -5131
rect 617 -5187 653 -5131
rect 525 -5349 653 -5187
rect 525 -5405 561 -5349
rect 617 -5405 653 -5349
rect 525 -5443 653 -5405
rect 305 -5995 881 -5955
rect 305 -6047 343 -5995
rect 395 -6047 791 -5995
rect 843 -6047 881 -5995
rect 305 -6213 881 -6047
rect 305 -6265 343 -6213
rect 395 -6265 791 -6213
rect 843 -6265 881 -6213
rect 305 -6306 881 -6265
rect 81 -7838 209 -7801
rect 81 -7894 117 -7838
rect 173 -7894 209 -7838
rect 81 -8056 209 -7894
rect 753 -7988 881 -6306
rect 81 -8112 117 -8056
rect 173 -8112 209 -8056
rect 81 -8274 209 -8112
rect 81 -8330 117 -8274
rect 173 -8330 209 -8274
rect 81 -8368 209 -8330
rect 81 -9797 209 -9760
rect 81 -9853 117 -9797
rect 173 -9853 209 -9797
rect 81 -10015 209 -9853
rect 81 -10071 117 -10015
rect 173 -10071 209 -10015
rect 81 -10233 209 -10071
rect 81 -10289 117 -10233
rect 173 -10289 209 -10233
rect 81 -10451 209 -10289
rect 81 -10507 117 -10451
rect 173 -10507 209 -10451
rect 81 -10545 209 -10507
<< via2 >>
rect 572 167 628 169
rect 572 115 574 167
rect 574 115 626 167
rect 626 115 628 167
rect 572 113 628 115
rect 572 -51 628 -49
rect 572 -103 574 -51
rect 574 -103 626 -51
rect 626 -103 628 -51
rect 572 -105 628 -103
rect 572 -269 628 -267
rect 572 -321 574 -269
rect 574 -321 626 -269
rect 626 -321 628 -269
rect 572 -323 628 -321
rect 572 -487 628 -485
rect 572 -539 574 -487
rect 574 -539 626 -487
rect 626 -539 628 -487
rect 572 -541 628 -539
rect 117 -2925 173 -2923
rect 117 -2977 119 -2925
rect 119 -2977 171 -2925
rect 171 -2977 173 -2925
rect 117 -2979 173 -2977
rect 117 -3143 173 -3141
rect 117 -3195 119 -3143
rect 119 -3195 171 -3143
rect 171 -3195 173 -3143
rect 117 -3197 173 -3195
rect 117 -3361 173 -3359
rect 117 -3413 119 -3361
rect 119 -3413 171 -3361
rect 171 -3413 173 -3361
rect 117 -3415 173 -3413
rect 565 -2925 621 -2923
rect 565 -2977 567 -2925
rect 567 -2977 619 -2925
rect 619 -2977 621 -2925
rect 565 -2979 621 -2977
rect 565 -3143 621 -3141
rect 565 -3195 567 -3143
rect 567 -3195 619 -3143
rect 619 -3195 621 -3143
rect 565 -3197 621 -3195
rect 565 -3361 621 -3359
rect 565 -3413 567 -3361
rect 567 -3413 619 -3361
rect 619 -3413 621 -3361
rect 565 -3415 621 -3413
rect 117 -4045 173 -4043
rect 117 -4097 119 -4045
rect 119 -4097 171 -4045
rect 171 -4097 173 -4045
rect 117 -4099 173 -4097
rect 117 -4263 173 -4261
rect 117 -4315 119 -4263
rect 119 -4315 171 -4263
rect 171 -4315 173 -4263
rect 117 -4317 173 -4315
rect 117 -4480 173 -4478
rect 117 -4532 119 -4480
rect 119 -4532 171 -4480
rect 171 -4532 173 -4480
rect 117 -4534 173 -4532
rect 117 -4698 173 -4696
rect 117 -4750 119 -4698
rect 119 -4750 171 -4698
rect 171 -4750 173 -4698
rect 117 -4752 173 -4750
rect 117 -4916 173 -4914
rect 117 -4968 119 -4916
rect 119 -4968 171 -4916
rect 171 -4968 173 -4916
rect 117 -4970 173 -4968
rect 117 -5133 173 -5131
rect 117 -5185 119 -5133
rect 119 -5185 171 -5133
rect 171 -5185 173 -5133
rect 117 -5187 173 -5185
rect 117 -5351 173 -5349
rect 117 -5403 119 -5351
rect 119 -5403 171 -5351
rect 171 -5403 173 -5351
rect 117 -5405 173 -5403
rect 561 -4045 617 -4043
rect 561 -4097 563 -4045
rect 563 -4097 615 -4045
rect 615 -4097 617 -4045
rect 561 -4099 617 -4097
rect 561 -4263 617 -4261
rect 561 -4315 563 -4263
rect 563 -4315 615 -4263
rect 615 -4315 617 -4263
rect 561 -4317 617 -4315
rect 561 -4480 617 -4478
rect 561 -4532 563 -4480
rect 563 -4532 615 -4480
rect 615 -4532 617 -4480
rect 561 -4534 617 -4532
rect 561 -4698 617 -4696
rect 561 -4750 563 -4698
rect 563 -4750 615 -4698
rect 615 -4750 617 -4698
rect 561 -4752 617 -4750
rect 561 -4916 617 -4914
rect 561 -4968 563 -4916
rect 563 -4968 615 -4916
rect 615 -4968 617 -4916
rect 561 -4970 617 -4968
rect 561 -5133 617 -5131
rect 561 -5185 563 -5133
rect 563 -5185 615 -5133
rect 615 -5185 617 -5133
rect 561 -5187 617 -5185
rect 561 -5351 617 -5349
rect 561 -5403 563 -5351
rect 563 -5403 615 -5351
rect 615 -5403 617 -5351
rect 561 -5405 617 -5403
rect 117 -7894 173 -7838
rect 117 -8112 173 -8056
rect 117 -8330 173 -8274
rect 117 -9853 173 -9797
rect 117 -10071 173 -10015
rect 117 -10289 173 -10233
rect 117 -10507 173 -10451
<< metal3 >>
rect -52 169 1106 327
rect -52 113 572 169
rect 628 113 1106 169
rect -52 -49 1106 113
rect -52 -105 572 -49
rect 628 -105 1106 -49
rect -52 -267 1106 -105
rect -52 -323 572 -267
rect 628 -323 1106 -267
rect -52 -485 1106 -323
rect -52 -541 572 -485
rect 628 -541 1106 -485
rect -52 -624 1106 -541
rect -58 -2923 1106 -2831
rect -58 -2979 117 -2923
rect 173 -2979 565 -2923
rect 621 -2979 1106 -2923
rect -58 -3141 1106 -2979
rect -58 -3197 117 -3141
rect 173 -3197 565 -3141
rect 621 -3197 1106 -3141
rect -58 -3359 1106 -3197
rect -58 -3415 117 -3359
rect 173 -3415 565 -3359
rect 621 -3415 1106 -3359
rect -58 -4043 1106 -3415
rect -58 -4099 117 -4043
rect 173 -4099 561 -4043
rect 617 -4099 1106 -4043
rect -58 -4261 1106 -4099
rect -58 -4317 117 -4261
rect 173 -4317 561 -4261
rect 617 -4317 1106 -4261
rect -58 -4478 1106 -4317
rect -58 -4534 117 -4478
rect 173 -4534 561 -4478
rect 617 -4534 1106 -4478
rect -58 -4696 1106 -4534
rect -58 -4752 117 -4696
rect 173 -4752 561 -4696
rect 617 -4752 1106 -4696
rect -58 -4914 1106 -4752
rect -58 -4970 117 -4914
rect 173 -4970 561 -4914
rect 617 -4970 1106 -4914
rect -58 -5131 1106 -4970
rect -58 -5187 117 -5131
rect 173 -5187 561 -5131
rect 617 -5187 1106 -5131
rect -58 -5349 1106 -5187
rect -58 -5405 117 -5349
rect 173 -5405 561 -5349
rect 617 -5405 1106 -5349
rect -58 -5553 1106 -5405
rect -1 -7838 963 -7728
rect -1 -7894 117 -7838
rect 173 -7894 963 -7838
rect -1 -8056 963 -7894
rect -1 -8112 117 -8056
rect 173 -8112 963 -8056
rect -1 -8274 963 -8112
rect -1 -8330 117 -8274
rect 173 -8330 963 -8274
rect -1 -8409 963 -8330
rect -67 -9797 1106 -9737
rect -67 -9853 117 -9797
rect 173 -9853 1106 -9797
rect -67 -10015 1106 -9853
rect -67 -10071 117 -10015
rect 173 -10071 1106 -10015
rect -67 -10233 1106 -10071
rect -67 -10289 117 -10233
rect 173 -10289 1106 -10233
rect -67 -10451 1106 -10289
rect -67 -10507 117 -10451
rect 173 -10507 1106 -10451
rect -67 -10645 1106 -10507
use M1_POLY24310589983261_64x8m81  M1_POLY24310589983261_64x8m81_0
timestamp 1666464484
transform 1 0 491 0 1 -3721
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_0
timestamp 1666464484
transform 1 0 817 0 1 -6130
box 0 0 1 1
use M2_M1$$43375660_64x8m81  M2_M1$$43375660_64x8m81_1
timestamp 1666464484
transform 1 0 369 0 1 -6130
box 0 0 1 1
use M2_M1$$43376684_64x8m81  M2_M1$$43376684_64x8m81_0
timestamp 1666464484
transform 1 0 817 0 1 -8524
box -63 -828 64 828
use M2_M1$$43379756_64x8m81  M2_M1$$43379756_64x8m81_0
timestamp 1666464484
transform 1 0 600 0 1 -186
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -3169
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_1
timestamp 1666464484
transform 1 0 593 0 1 -3169
box 0 0 1 1
use M2_M1$$43380780_64x8m81  M2_M1$$43380780_64x8m81_2
timestamp 1666464484
transform 1 0 367 0 1 -428
box 0 0 1 1
use M2_M1$$47327276_64x8m81  M2_M1$$47327276_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -9172
box -65 -1373 65 1373
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -4724
box 0 0 1 1
use M2_M1$$47515692_64x8m81  M2_M1$$47515692_64x8m81_1
timestamp 1666464484
transform 1 0 589 0 1 -4724
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -3169
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_1
timestamp 1666464484
transform 1 0 593 0 1 -3169
box 0 0 1 1
use M3_M2$$47108140_64x8m81  M3_M2$$47108140_64x8m81_2
timestamp 1666464484
transform 1 0 145 0 1 -8084
box 0 0 1 1
use M3_M2$$47332396_64x8m81  M3_M2$$47332396_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -4724
box 0 0 1 1
use M3_M2$$47332396_64x8m81  M3_M2$$47332396_64x8m81_1
timestamp 1666464484
transform 1 0 589 0 1 -4724
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_0
timestamp 1666464484
transform 1 0 145 0 1 -10152
box 0 0 1 1
use M3_M2$$47333420_64x8m81  M3_M2$$47333420_64x8m81_1
timestamp 1666464484
transform 1 0 600 0 1 -186
box 0 0 1 1
use nmos_1p2$$47514668_64x8m81  nmos_1p2$$47514668_64x8m81_0
timestamp 1666464484
transform 1 0 228 0 -1 -136
box -119 -73 177 980
use nmos_1p2$$47514668_64x8m81  nmos_1p2$$47514668_64x8m81_1
timestamp 1666464484
transform 1 0 452 0 -1 -136
box -119 -73 177 980
use nmos_1p2$$47514668_64x8m81  nmos_1p2$$47514668_64x8m81_2
timestamp 1666464484
transform 1 0 676 0 -1 -136
box -119 -73 177 980
use pmos_1p2$$47512620_64x8m81  pmos_1p2$$47512620_64x8m81_0
timestamp 1666464484
transform 1 0 676 0 1 -6314
box -286 -142 344 2227
use pmos_1p2$$47512620_64x8m81  pmos_1p2$$47512620_64x8m81_1
timestamp 1666464484
transform 1 0 452 0 1 -6314
box -286 -142 344 2227
use pmos_1p2$$47512620_64x8m81  pmos_1p2$$47512620_64x8m81_2
timestamp 1666464484
transform 1 0 228 0 1 -6314
box -286 -142 344 2227
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_0
timestamp 1666464484
transform 1 0 452 0 -1 -1324
box -286 -141 344 2409
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_1
timestamp 1666464484
transform 1 0 676 0 -1 -1324
box -286 -141 344 2409
use pmos_1p2$$47513644_64x8m81  pmos_1p2$$47513644_64x8m81_2
timestamp 1666464484
transform 1 0 228 0 -1 -1324
box -286 -141 344 2409
<< properties >>
string GDS_END 479422
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 472814
<< end >>
