magic
tech gf180mcuB
timestamp 1666464484
<< metal1 >>
rect 0 111 102 123
rect 11 70 16 111
rect 11 57 21 63
rect 45 51 50 104
rect 62 91 67 104
rect 62 81 68 91
rect 45 43 57 51
rect 11 12 16 36
rect 45 19 50 43
rect 62 19 67 81
rect 85 51 90 104
rect 85 43 95 51
rect 85 19 90 43
rect 0 0 102 12
<< obsm1 >>
rect 28 67 33 104
rect 28 61 39 67
rect 28 46 33 61
rect 28 40 40 46
rect 28 19 33 40
rect 73 58 79 69
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 60 82 70 90
rect 11 56 21 64
rect 47 43 57 51
rect 85 43 95 51
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
<< obsm2 >>
rect 29 67 39 68
rect 71 67 81 68
rect 29 61 81 67
rect 29 60 39 61
rect 71 60 81 61
<< labels >>
rlabel metal2 s 47 43 57 51 6 A
port 1 nsew signal input
rlabel metal1 s 45 19 50 104 6 A
port 1 nsew signal input
rlabel metal1 s 45 43 57 51 6 A
port 1 nsew signal input
rlabel metal2 s 85 43 95 51 6 B
port 2 nsew signal input
rlabel metal1 s 85 19 90 104 6 B
port 2 nsew signal input
rlabel metal1 s 85 43 95 51 6 B
port 2 nsew signal input
rlabel metal2 s 11 56 21 64 6 Sel
port 3 nsew signal output
rlabel metal1 s 11 57 21 63 6 Sel
port 3 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 11 70 16 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 111 102 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 11 0 16 36 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 102 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 60 82 70 90 6 Y
port 6 nsew signal output
rlabel metal1 s 62 19 67 104 6 Y
port 6 nsew signal output
rlabel metal1 s 62 81 68 91 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 102 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
