magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 4816 844
rect 69 536 115 622
rect 486 618 554 724
rect 945 536 991 622
rect 1382 618 1450 724
rect 1841 536 1887 622
rect 2005 536 2051 622
rect 2198 618 2266 724
rect 2433 536 2479 622
rect 2646 618 2714 724
rect 3318 657 3386 724
rect 3447 611 4147 662
rect 4214 657 4282 724
rect 2870 582 4756 611
rect 2870 565 3493 582
rect 4101 565 4756 582
rect 2870 536 2938 565
rect 69 472 2938 536
rect 3594 519 4022 536
rect 124 360 318 424
rect 368 360 1542 424
rect 270 314 318 360
rect 1588 354 1894 424
rect 2023 360 2832 424
rect 1588 314 1634 354
rect 270 268 1634 314
rect 2881 244 2938 472
rect 3003 473 4022 519
rect 3003 320 3049 473
rect 3143 360 3585 424
rect 3664 382 3732 473
rect 3868 428 4022 473
rect 3868 382 4684 428
rect 3535 336 3585 360
rect 4477 358 4684 382
rect 3535 290 4376 336
rect 2881 198 4506 244
rect 4612 224 4684 358
rect 38 60 106 127
rect 485 60 554 127
rect 933 60 1002 127
rect 1381 60 1450 127
rect 1829 60 1898 127
rect 0 -60 4816 60
<< obsm1 >>
rect 1757 219 2714 244
rect 244 198 2714 219
rect 244 173 1807 198
rect 1972 106 4776 152
<< labels >>
rlabel metal1 s 3594 519 4022 536 6 A1
port 1 nsew default input
rlabel metal1 s 3003 473 4022 519 6 A1
port 1 nsew default input
rlabel metal1 s 3868 428 4022 473 6 A1
port 1 nsew default input
rlabel metal1 s 3664 428 3732 473 6 A1
port 1 nsew default input
rlabel metal1 s 3003 428 3049 473 6 A1
port 1 nsew default input
rlabel metal1 s 3868 382 4684 428 6 A1
port 1 nsew default input
rlabel metal1 s 3664 382 3732 428 6 A1
port 1 nsew default input
rlabel metal1 s 3003 382 3049 428 6 A1
port 1 nsew default input
rlabel metal1 s 4477 358 4684 382 6 A1
port 1 nsew default input
rlabel metal1 s 3003 358 3049 382 6 A1
port 1 nsew default input
rlabel metal1 s 4612 320 4684 358 6 A1
port 1 nsew default input
rlabel metal1 s 3003 320 3049 358 6 A1
port 1 nsew default input
rlabel metal1 s 4612 224 4684 320 6 A1
port 1 nsew default input
rlabel metal1 s 3143 360 3585 424 6 A2
port 2 nsew default input
rlabel metal1 s 3535 336 3585 360 6 A2
port 2 nsew default input
rlabel metal1 s 3535 290 4376 336 6 A2
port 2 nsew default input
rlabel metal1 s 1588 360 1894 424 6 B1
port 3 nsew default input
rlabel metal1 s 124 360 318 424 6 B1
port 3 nsew default input
rlabel metal1 s 1588 354 1894 360 6 B1
port 3 nsew default input
rlabel metal1 s 270 354 318 360 6 B1
port 3 nsew default input
rlabel metal1 s 1588 314 1634 354 6 B1
port 3 nsew default input
rlabel metal1 s 270 314 318 354 6 B1
port 3 nsew default input
rlabel metal1 s 270 268 1634 314 6 B1
port 3 nsew default input
rlabel metal1 s 368 360 1542 424 6 B2
port 4 nsew default input
rlabel metal1 s 2023 360 2832 424 6 C
port 5 nsew default input
rlabel metal1 s 3447 622 4147 662 6 ZN
port 6 nsew default output
rlabel metal1 s 3447 611 4147 622 6 ZN
port 6 nsew default output
rlabel metal1 s 2433 611 2479 622 6 ZN
port 6 nsew default output
rlabel metal1 s 2005 611 2051 622 6 ZN
port 6 nsew default output
rlabel metal1 s 1841 611 1887 622 6 ZN
port 6 nsew default output
rlabel metal1 s 945 611 991 622 6 ZN
port 6 nsew default output
rlabel metal1 s 69 611 115 622 6 ZN
port 6 nsew default output
rlabel metal1 s 2870 582 4756 611 6 ZN
port 6 nsew default output
rlabel metal1 s 2433 582 2479 611 6 ZN
port 6 nsew default output
rlabel metal1 s 2005 582 2051 611 6 ZN
port 6 nsew default output
rlabel metal1 s 1841 582 1887 611 6 ZN
port 6 nsew default output
rlabel metal1 s 945 582 991 611 6 ZN
port 6 nsew default output
rlabel metal1 s 69 582 115 611 6 ZN
port 6 nsew default output
rlabel metal1 s 4101 565 4756 582 6 ZN
port 6 nsew default output
rlabel metal1 s 2870 565 3493 582 6 ZN
port 6 nsew default output
rlabel metal1 s 2433 565 2479 582 6 ZN
port 6 nsew default output
rlabel metal1 s 2005 565 2051 582 6 ZN
port 6 nsew default output
rlabel metal1 s 1841 565 1887 582 6 ZN
port 6 nsew default output
rlabel metal1 s 945 565 991 582 6 ZN
port 6 nsew default output
rlabel metal1 s 69 565 115 582 6 ZN
port 6 nsew default output
rlabel metal1 s 2870 536 2938 565 6 ZN
port 6 nsew default output
rlabel metal1 s 2433 536 2479 565 6 ZN
port 6 nsew default output
rlabel metal1 s 2005 536 2051 565 6 ZN
port 6 nsew default output
rlabel metal1 s 1841 536 1887 565 6 ZN
port 6 nsew default output
rlabel metal1 s 945 536 991 565 6 ZN
port 6 nsew default output
rlabel metal1 s 69 536 115 565 6 ZN
port 6 nsew default output
rlabel metal1 s 69 472 2938 536 6 ZN
port 6 nsew default output
rlabel metal1 s 2881 244 2938 472 6 ZN
port 6 nsew default output
rlabel metal1 s 2881 198 4506 244 6 ZN
port 6 nsew default output
rlabel metal1 s 0 724 4816 844 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4214 657 4282 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3318 657 3386 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2646 657 2714 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2198 657 2266 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1382 657 1450 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 486 657 554 724 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2646 618 2714 657 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2198 618 2266 657 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1382 618 1450 657 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 486 618 554 657 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1829 60 1898 127 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1381 60 1450 127 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 933 60 1002 127 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 485 60 554 127 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 38 60 106 127 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 4816 60 8 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 4816 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 120256
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 112020
<< end >>
