magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -169 463 170 502
rect -169 407 -134 463
rect -78 407 78 463
rect 134 407 170 463
rect -169 246 170 407
rect -169 190 -134 246
rect -78 190 78 246
rect 134 190 170 246
rect -169 28 170 190
rect -169 -28 -134 28
rect -78 -28 78 28
rect 134 -28 170 28
rect -169 -190 170 -28
rect -169 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 170 -190
rect -169 -407 170 -246
rect -169 -463 -134 -407
rect -78 -463 78 -407
rect 134 -463 170 -407
rect -169 -502 170 -463
<< via2 >>
rect -134 407 -78 463
rect 78 407 134 463
rect -134 190 -78 246
rect 78 190 134 246
rect -134 -28 -78 28
rect 78 -28 134 28
rect -134 -246 -78 -190
rect 78 -246 134 -190
rect -134 -463 -78 -407
rect 78 -463 134 -407
<< metal3 >>
rect -170 463 170 502
rect -170 407 -134 463
rect -78 407 78 463
rect 134 407 170 463
rect -170 246 170 407
rect -170 190 -134 246
rect -78 190 78 246
rect 134 190 170 246
rect -170 28 170 190
rect -170 -28 -134 28
rect -78 -28 78 28
rect 134 -28 170 28
rect -170 -190 170 -28
rect -170 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 170 -190
rect -170 -407 170 -246
rect -170 -463 -134 -407
rect -78 -463 78 -407
rect 134 -463 170 -407
rect -170 -502 170 -463
<< properties >>
string GDS_END 1112604
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1111832
<< end >>
