magic
tech gf180mcuC
timestamp 1667403419
<< metal1 >>
rect 0 111 190 123
rect 29 86 34 111
rect 107 75 112 111
rect 37 57 47 63
rect 68 57 78 66
rect 114 60 124 66
rect 29 12 37 30
rect 156 84 161 111
rect 104 12 112 29
rect 173 64 178 104
rect 173 63 181 64
rect 173 57 183 63
rect 173 56 181 57
rect 156 12 161 29
rect 173 19 178 56
rect 0 0 190 12
<< obsm1 >>
rect 12 51 17 104
rect 63 81 68 104
rect 23 76 68 81
rect 23 66 28 76
rect 124 78 129 104
rect 124 73 134 78
rect 22 60 31 66
rect 10 50 17 51
rect 7 44 17 50
rect 9 43 17 44
rect 12 19 17 43
rect 23 43 28 60
rect 52 60 62 66
rect 54 52 60 60
rect 83 52 93 55
rect 54 49 93 52
rect 54 47 91 49
rect 100 47 110 53
rect 54 46 90 47
rect 23 38 48 43
rect 43 29 48 38
rect 84 39 90 46
rect 129 45 134 73
rect 139 72 144 104
rect 139 67 166 72
rect 144 47 154 53
rect 124 40 134 45
rect 160 42 166 67
rect 124 39 129 40
rect 84 34 129 39
rect 63 29 68 31
rect 43 24 68 29
rect 63 19 68 24
rect 124 19 129 34
rect 139 37 166 42
rect 139 19 144 37
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 82 118 90 119
rect 106 118 114 119
rect 130 118 138 119
rect 154 118 162 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 81 112 91 118
rect 105 112 115 118
rect 129 112 139 118
rect 153 112 163 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 82 111 90 112
rect 106 111 114 112
rect 130 111 138 112
rect 154 111 162 112
rect 114 66 124 67
rect 70 64 124 66
rect 37 56 47 64
rect 69 63 124 64
rect 174 63 182 64
rect 68 60 124 63
rect 68 57 78 60
rect 114 59 124 60
rect 173 57 183 63
rect 69 56 77 57
rect 174 56 182 57
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
<< obsm2 >>
rect 101 53 109 54
rect 144 53 154 54
rect 7 50 17 51
rect 92 50 154 53
rect 7 47 154 50
rect 7 46 109 47
rect 144 46 154 47
rect 7 44 98 46
rect 7 43 17 44
<< labels >>
rlabel metal2 s 69 56 77 64 6 CLKN
port 1 nsew clock input
rlabel metal2 s 68 57 78 63 6 CLKN
port 1 nsew clock input
rlabel metal2 s 70 60 124 66 6 CLKN
port 1 nsew clock input
rlabel metal2 s 114 59 124 67 6 CLKN
port 1 nsew clock input
rlabel metal1 s 68 57 78 66 6 CLKN
port 1 nsew clock input
rlabel metal1 s 114 60 124 66 6 CLKN
port 1 nsew clock input
rlabel metal2 s 37 56 47 64 6 D
port 2 nsew signal input
rlabel metal1 s 37 57 47 63 6 D
port 2 nsew signal input
rlabel metal2 s 174 56 182 64 6 Q
port 3 nsew signal output
rlabel metal2 s 173 57 183 63 6 Q
port 3 nsew signal output
rlabel metal1 s 173 19 178 104 6 Q
port 3 nsew signal output
rlabel metal1 s 173 56 181 64 6 Q
port 3 nsew signal output
rlabel metal1 s 173 57 183 63 6 Q
port 3 nsew signal output
rlabel metal2 s 10 111 18 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 82 111 90 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 81 112 91 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 106 111 114 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 105 112 115 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 130 111 138 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 129 112 139 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 154 111 162 119 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 153 112 163 118 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 29 86 34 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 107 75 112 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 156 84 161 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 111 190 123 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 29 0 37 30 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 104 0 112 29 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 156 0 161 29 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 0 0 190 12 6 VSS
port 5 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 190 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
