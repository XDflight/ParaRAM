magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -78 23 1817 80
rect -78 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1817 23
rect -78 -80 1817 -23
<< psubdiffcont >>
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect 1242 -23 1288 23
rect 1400 -23 1446 23
rect 1558 -23 1604 23
rect 1716 -23 1762 23
<< metal1 >>
rect -58 23 1797 60
rect -58 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1242 23
rect 1288 -23 1400 23
rect 1446 -23 1558 23
rect 1604 -23 1716 23
rect 1762 -23 1797 23
rect -58 -60 1797 -23
<< properties >>
string GDS_END 2526670
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2525706
<< end >>
