magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -1386 156 -1226 157
rect -1386 102 1386 156
rect -1386 56 -1329 102
rect -1283 56 -1166 102
rect -1120 56 -1003 102
rect -957 56 -839 102
rect -793 56 -676 102
rect -630 56 -513 102
rect -467 56 -350 102
rect -304 56 -186 102
rect -140 56 -23 102
rect 23 56 140 102
rect 186 56 304 102
rect 350 56 467 102
rect 513 56 630 102
rect 676 56 793 102
rect 839 56 957 102
rect 1003 56 1120 102
rect 1166 56 1283 102
rect 1329 56 1386 102
rect -1386 -56 1386 56
rect -1386 -102 -1329 -56
rect -1283 -102 -1166 -56
rect -1120 -102 -1003 -56
rect -957 -102 -839 -56
rect -793 -102 -676 -56
rect -630 -102 -513 -56
rect -467 -102 -350 -56
rect -304 -102 -186 -56
rect -140 -102 -23 -56
rect 23 -102 140 -56
rect 186 -102 304 -56
rect 350 -102 467 -56
rect 513 -102 630 -56
rect 676 -102 793 -56
rect 839 -102 957 -56
rect 1003 -102 1120 -56
rect 1166 -102 1283 -56
rect 1329 -102 1386 -56
rect -1386 -157 1386 -102
<< psubdiffcont >>
rect -1329 56 -1283 102
rect -1166 56 -1120 102
rect -1003 56 -957 102
rect -839 56 -793 102
rect -676 56 -630 102
rect -513 56 -467 102
rect -350 56 -304 102
rect -186 56 -140 102
rect -23 56 23 102
rect 140 56 186 102
rect 304 56 350 102
rect 467 56 513 102
rect 630 56 676 102
rect 793 56 839 102
rect 957 56 1003 102
rect 1120 56 1166 102
rect 1283 56 1329 102
rect -1329 -102 -1283 -56
rect -1166 -102 -1120 -56
rect -1003 -102 -957 -56
rect -839 -102 -793 -56
rect -676 -102 -630 -56
rect -513 -102 -467 -56
rect -350 -102 -304 -56
rect -186 -102 -140 -56
rect -23 -102 23 -56
rect 140 -102 186 -56
rect 304 -102 350 -56
rect 467 -102 513 -56
rect 630 -102 676 -56
rect 793 -102 839 -56
rect 957 -102 1003 -56
rect 1120 -102 1166 -56
rect 1283 -102 1329 -56
<< metal1 >>
rect -1366 102 1366 137
rect -1366 56 -1329 102
rect -1283 56 -1166 102
rect -1120 56 -1003 102
rect -957 56 -839 102
rect -793 56 -676 102
rect -630 56 -513 102
rect -467 56 -350 102
rect -304 56 -186 102
rect -140 56 -23 102
rect 23 56 140 102
rect 186 56 304 102
rect 350 56 467 102
rect 513 56 630 102
rect 676 56 793 102
rect 839 56 957 102
rect 1003 56 1120 102
rect 1166 56 1283 102
rect 1329 56 1366 102
rect -1366 -56 1366 56
rect -1366 -102 -1329 -56
rect -1283 -102 -1166 -56
rect -1120 -102 -1003 -56
rect -957 -102 -839 -56
rect -793 -102 -676 -56
rect -630 -102 -513 -56
rect -467 -102 -350 -56
rect -304 -102 -186 -56
rect -140 -102 -23 -56
rect 23 -102 140 -56
rect 186 -102 304 -56
rect 350 -102 467 -56
rect 513 -102 630 -56
rect 676 -102 793 -56
rect 839 -102 957 -56
rect 1003 -102 1120 -56
rect 1166 -102 1283 -56
rect 1329 -102 1366 -56
rect -1366 -137 1366 -102
<< properties >>
string GDS_END 809512
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 807092
<< end >>
