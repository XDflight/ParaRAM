magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -143 106 143 112
rect -143 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 143 106
rect -143 44 143 80
rect -143 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 143 44
rect -143 -18 143 18
rect -143 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 143 -18
rect -143 -80 143 -44
rect -143 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 143 -80
rect -143 -112 143 -106
<< via1 >>
rect -137 80 -111 106
rect -75 80 -49 106
rect -13 80 13 106
rect 49 80 75 106
rect 111 80 137 106
rect -137 18 -111 44
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect 111 18 137 44
rect -137 -44 -111 -18
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect 111 -44 137 -18
rect -137 -106 -111 -80
rect -75 -106 -49 -80
rect -13 -106 13 -80
rect 49 -106 75 -80
rect 111 -106 137 -80
<< metal2 >>
rect -143 106 143 112
rect -143 80 -137 106
rect -111 80 -75 106
rect -49 80 -13 106
rect 13 80 49 106
rect 75 80 111 106
rect 137 80 143 106
rect -143 44 143 80
rect -143 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 143 44
rect -143 -18 143 18
rect -143 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 143 -18
rect -143 -80 143 -44
rect -143 -106 -137 -80
rect -111 -106 -75 -80
rect -49 -106 -13 -80
rect 13 -106 49 -80
rect 75 -106 111 -80
rect 137 -106 143 -80
rect -143 -112 143 -106
<< properties >>
string GDS_END 2650976
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2649564
<< end >>
