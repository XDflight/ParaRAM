magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal3 >>
rect -511 630 489 2430
rect 714 1822 1714 2430
use M2_M14310591302017_512x8m81  M2_M14310591302017_512x8m81_0
timestamp 1666464484
transform 1 0 1214 0 1 1986
box -472 -162 472 162
use M3_M24310591302016_512x8m81  M3_M24310591302016_512x8m81_0
timestamp 1666464484
transform 1 0 1214 0 1 1986
box -472 -162 472 162
use M3_M24310591302042_512x8m81  M3_M24310591302042_512x8m81_0
timestamp 1666464484
transform 1 0 -12 0 1 1126
box -472 -472 472 472
<< properties >>
string GDS_END 2876104
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2875836
string path -0.055 3.150 -0.055 12.150 
<< end >>
