magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 784 844
rect 76 506 122 724
rect 280 556 326 676
rect 473 626 541 724
rect 676 556 734 676
rect 280 472 734 556
rect 24 352 213 430
rect 132 211 213 352
rect 76 60 122 161
rect 356 110 428 392
rect 580 110 642 392
rect 688 131 734 472
rect 0 -60 784 60
<< labels >>
rlabel metal1 s 580 110 642 392 6 A1
port 1 nsew default input
rlabel metal1 s 356 110 428 392 6 A2
port 2 nsew default input
rlabel metal1 s 24 352 213 430 6 A3
port 3 nsew default input
rlabel metal1 s 132 211 213 352 6 A3
port 3 nsew default input
rlabel metal1 s 676 556 734 676 6 ZN
port 4 nsew default output
rlabel metal1 s 280 556 326 676 6 ZN
port 4 nsew default output
rlabel metal1 s 280 472 734 556 6 ZN
port 4 nsew default output
rlabel metal1 s 688 131 734 472 6 ZN
port 4 nsew default output
rlabel metal1 s 0 724 784 844 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 473 626 541 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 76 626 122 724 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 76 506 122 626 6 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 76 60 122 161 6 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 784 60 8 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 784 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 698848
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 696016
<< end >>
