magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 918 896 1098
rect 253 710 299 918
rect 30 466 194 542
rect 126 400 194 466
rect 497 603 543 872
rect 701 710 747 918
rect 497 546 656 603
rect 596 318 656 546
rect 466 242 656 318
rect 273 90 319 233
rect 466 142 543 242
rect 721 90 767 304
rect 0 -90 896 90
<< obsm1 >>
rect 49 664 95 872
rect 49 618 286 664
rect 240 500 286 618
rect 240 454 550 500
rect 240 325 286 454
rect 49 279 286 325
rect 49 142 95 279
<< labels >>
rlabel metal1 s 30 466 194 542 6 I
port 1 nsew default input
rlabel metal1 s 126 400 194 466 6 I
port 1 nsew default input
rlabel metal1 s 497 603 543 872 6 Z
port 2 nsew default output
rlabel metal1 s 497 546 656 603 6 Z
port 2 nsew default output
rlabel metal1 s 596 318 656 546 6 Z
port 2 nsew default output
rlabel metal1 s 466 242 656 318 6 Z
port 2 nsew default output
rlabel metal1 s 466 142 543 242 6 Z
port 2 nsew default output
rlabel metal1 s 0 918 896 1098 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 701 710 747 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 253 710 299 918 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 721 233 767 304 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 721 90 767 233 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 233 6 VSS
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 896 90 8 VSS
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 896 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1240604
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 1237222
<< end >>
