magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 6583 14608 9560 15532
rect 13849 15258 15116 15548
rect 13849 15181 15441 15258
rect 10186 14617 10786 14689
rect 13850 14608 15441 15181
rect 6583 14558 8962 14608
rect 16520 14576 21087 15503
<< mvndiff >>
rect 2123 14460 2278 14848
rect 25490 14460 25646 14848
<< mvpsubdiff >>
rect 15782 15382 16254 15439
rect 15782 15336 15837 15382
rect 15883 15336 15995 15382
rect 16041 15336 16153 15382
rect 16199 15336 16254 15382
rect 15782 15279 16254 15336
<< mvnsubdiff >>
rect 13985 15382 14931 15439
rect 13985 15336 14040 15382
rect 14086 15336 14198 15382
rect 14244 15336 14356 15382
rect 14402 15336 14514 15382
rect 14560 15336 14673 15382
rect 14719 15336 14831 15382
rect 14877 15336 14931 15382
rect 13985 15279 14931 15336
<< mvpsubdiffcont >>
rect 15837 15336 15883 15382
rect 15995 15336 16041 15382
rect 16153 15336 16199 15382
<< mvnsubdiffcont >>
rect 14040 15336 14086 15382
rect 14198 15336 14244 15382
rect 14356 15336 14402 15382
rect 14514 15336 14560 15382
rect 14673 15336 14719 15382
rect 14831 15336 14877 15382
<< polysilicon >>
rect 13623 15316 13801 15335
rect 13623 15270 13642 15316
rect 13782 15270 13801 15316
rect 15364 15364 15467 15383
rect 15364 15318 15390 15364
rect 15436 15318 15467 15364
rect 13623 15251 13801 15270
rect 6556 15096 6690 15216
rect 9314 15118 9448 15223
rect 6556 14992 6659 15096
rect 6374 14872 6690 14992
rect 9314 14978 9358 15118
rect 9404 14978 9448 15118
rect 11998 15031 12082 15050
rect 11998 14992 12017 15031
rect 9314 14873 9448 14978
rect 11043 14872 11385 14992
rect 11914 14891 12017 14992
rect 12063 14891 12082 15031
rect 11914 14872 12082 14891
rect 13664 14873 13768 15251
rect 15364 14992 15467 15318
rect 18271 15106 18355 15216
rect 13915 14872 13986 14992
rect 15305 14872 15467 14992
rect 15583 15071 15667 15090
rect 15583 14931 15602 15071
rect 15648 14992 15667 15071
rect 15648 14931 15755 14992
rect 15583 14872 15755 14931
rect 16255 14872 16656 14992
rect 17975 14872 18045 14992
rect 18271 14966 18290 15106
rect 18336 14966 18355 15106
rect 18271 14872 18355 14966
rect 21010 14992 21113 15216
rect 21010 14872 21325 14992
rect 23347 14872 23417 14992
<< polycontact >>
rect 13642 15270 13782 15316
rect 15390 15318 15436 15364
rect 9358 14978 9404 15118
rect 12017 14891 12063 15031
rect 15602 14931 15648 15071
rect 18290 14966 18336 15106
<< metal1 >>
rect 2123 14716 4017 15367
rect 4324 15052 6336 15439
rect 6728 15306 7700 15346
rect 6728 15254 6766 15306
rect 6818 15254 6977 15306
rect 7029 15254 7188 15306
rect 7240 15254 7399 15306
rect 7451 15254 7610 15306
rect 7662 15254 7700 15306
rect 6728 15214 7700 15254
rect 11385 15331 11913 15419
rect 11385 15279 11575 15331
rect 11627 15279 11755 15331
rect 11807 15279 11913 15331
rect 9323 15118 9439 15185
rect 6482 14988 6767 15108
rect 4335 14845 5307 14885
rect 6482 14877 6598 14988
rect 9323 14978 9358 15118
rect 9404 14978 9439 15118
rect 10338 15108 10888 15115
rect 10337 15074 10888 15108
rect 10337 15022 10376 15074
rect 10428 15022 10587 15074
rect 10639 15022 10798 15074
rect 10850 15022 10888 15074
rect 10337 14988 10888 15022
rect 11385 15113 11913 15279
rect 13531 15382 14912 15419
rect 15755 15418 16283 15419
rect 13531 15378 14040 15382
rect 13531 15326 14033 15378
rect 14086 15336 14198 15382
rect 14244 15378 14356 15382
rect 14085 15326 14244 15336
rect 14296 15336 14356 15378
rect 14402 15378 14514 15382
rect 14402 15336 14455 15378
rect 14296 15326 14455 15336
rect 14507 15336 14514 15378
rect 14560 15336 14673 15382
rect 14719 15336 14831 15382
rect 14877 15336 14912 15382
rect 14507 15326 14912 15336
rect 13531 15317 14912 15326
rect 13531 15265 13569 15317
rect 13621 15316 13781 15317
rect 13621 15270 13642 15316
rect 13833 15299 14912 15317
rect 15061 15382 16283 15418
rect 15061 15378 15837 15382
rect 15061 15326 15100 15378
rect 15152 15326 15311 15378
rect 15363 15364 15522 15378
rect 15363 15326 15390 15364
rect 15061 15318 15390 15326
rect 15436 15326 15522 15364
rect 15574 15326 15733 15378
rect 15785 15336 15837 15378
rect 15883 15336 15995 15382
rect 16041 15336 16153 15382
rect 16199 15336 16283 15382
rect 20112 15340 20874 15346
rect 15785 15326 16283 15336
rect 15436 15318 16283 15326
rect 13833 15286 14545 15299
rect 13833 15285 14040 15286
rect 15061 15285 16283 15318
rect 13621 15265 13781 15270
rect 13833 15265 13871 15285
rect 13531 15224 13871 15265
rect 11385 15061 11575 15113
rect 11627 15061 11755 15113
rect 11807 15061 11913 15113
rect 15591 15071 15659 15082
rect 11385 15021 11913 15061
rect 12006 15031 12334 15068
rect 10338 14982 10888 14988
rect 4335 14793 4373 14845
rect 4425 14793 4584 14845
rect 4636 14793 4795 14845
rect 4847 14793 5006 14845
rect 5058 14793 5217 14845
rect 5269 14793 5307 14845
rect 4335 14753 5307 14793
rect 6240 14757 6598 14877
rect 6728 14843 7700 14883
rect 6728 14791 6766 14843
rect 6818 14791 6977 14843
rect 7029 14791 7188 14843
rect 7240 14791 7399 14843
rect 7451 14791 7610 14843
rect 7662 14791 7700 14843
rect 6728 14751 7700 14791
rect 9323 14877 9439 14978
rect 12006 14891 12017 15031
rect 12063 15022 12334 15031
rect 13509 15022 14174 15068
rect 15591 15067 15602 15071
rect 12063 14891 12074 15022
rect 15268 15021 15602 15067
rect 15591 14931 15602 15021
rect 15648 14931 15659 15071
rect 15755 14988 16283 15285
rect 16656 15306 20942 15340
rect 16656 15254 20151 15306
rect 20203 15254 20362 15306
rect 20414 15254 20573 15306
rect 20625 15254 20784 15306
rect 20836 15254 20942 15306
rect 16656 15220 20942 15254
rect 16656 15036 17974 15220
rect 20112 15213 20874 15220
rect 18279 15106 18347 15117
rect 15591 14920 15659 14931
rect 18279 14966 18290 15106
rect 18336 14966 18347 15106
rect 20898 15021 21184 15067
rect 18279 14955 18347 14966
rect 12006 14880 12074 14891
rect 9323 14757 11913 14877
rect 12294 14843 13478 14884
rect 18279 14877 18346 14955
rect 12294 14791 12333 14843
rect 12385 14791 12544 14843
rect 12596 14791 12755 14843
rect 12807 14791 12966 14843
rect 13018 14791 13177 14843
rect 13229 14791 13387 14843
rect 13439 14791 13478 14843
rect 13570 14798 14174 14844
rect 12294 14750 13478 14791
rect 15755 14757 18346 14877
rect 20112 14843 20874 14883
rect 20112 14791 20151 14843
rect 20203 14791 20362 14843
rect 20414 14791 20573 14843
rect 20625 14791 20784 14843
rect 20836 14791 20874 14843
rect 21067 14843 21184 15021
rect 21324 15002 23346 15419
rect 22366 14843 23338 14883
rect 21067 14797 21425 14843
rect 20112 14750 20874 14791
rect 22366 14791 22404 14843
rect 22456 14791 22615 14843
rect 22667 14791 22826 14843
rect 22878 14791 23037 14843
rect 23089 14791 23248 14843
rect 23300 14791 23338 14843
rect 22366 14751 23338 14791
rect 23751 14716 25646 15367
rect 2123 14465 2278 14716
rect 25490 14465 25646 14716
<< via1 >>
rect 6766 15254 6818 15306
rect 6977 15254 7029 15306
rect 7188 15254 7240 15306
rect 7399 15254 7451 15306
rect 7610 15254 7662 15306
rect 11575 15279 11627 15331
rect 11755 15279 11807 15331
rect 10376 15022 10428 15074
rect 10587 15022 10639 15074
rect 10798 15022 10850 15074
rect 14033 15336 14040 15378
rect 14040 15336 14085 15378
rect 14033 15326 14085 15336
rect 14244 15326 14296 15378
rect 14455 15326 14507 15378
rect 13569 15265 13621 15317
rect 13781 15316 13833 15317
rect 13781 15270 13782 15316
rect 13782 15270 13833 15316
rect 15100 15326 15152 15378
rect 15311 15326 15363 15378
rect 15522 15326 15574 15378
rect 15733 15326 15785 15378
rect 13781 15265 13833 15270
rect 11575 15061 11627 15113
rect 11755 15061 11807 15113
rect 4373 14793 4425 14845
rect 4584 14793 4636 14845
rect 4795 14793 4847 14845
rect 5006 14793 5058 14845
rect 5217 14793 5269 14845
rect 6766 14791 6818 14843
rect 6977 14791 7029 14843
rect 7188 14791 7240 14843
rect 7399 14791 7451 14843
rect 7610 14791 7662 14843
rect 20151 15254 20203 15306
rect 20362 15254 20414 15306
rect 20573 15254 20625 15306
rect 20784 15254 20836 15306
rect 12333 14791 12385 14843
rect 12544 14791 12596 14843
rect 12755 14791 12807 14843
rect 12966 14791 13018 14843
rect 13177 14791 13229 14843
rect 13387 14791 13439 14843
rect 20151 14791 20203 14843
rect 20362 14791 20414 14843
rect 20573 14791 20625 14843
rect 20784 14791 20836 14843
rect 22404 14791 22456 14843
rect 22615 14791 22667 14843
rect 22826 14791 22878 14843
rect 23037 14791 23089 14843
rect 23248 14791 23300 14843
<< metal2 >>
rect 2092 14413 4211 15476
rect 5550 15328 6347 15401
rect 5550 15272 5611 15328
rect 5667 15272 5822 15328
rect 5878 15272 6033 15328
rect 6089 15272 6244 15328
rect 6300 15272 6347 15328
rect 4334 14847 5307 14886
rect 4334 14791 4371 14847
rect 4427 14791 4582 14847
rect 4638 14791 4793 14847
rect 4849 14791 5004 14847
rect 5060 14791 5215 14847
rect 5271 14791 5307 14847
rect 4334 14753 5307 14791
rect 5550 14413 6347 15272
rect 6451 15306 7738 15401
rect 6451 15254 6766 15306
rect 6818 15254 6977 15306
rect 7029 15254 7188 15306
rect 7240 15254 7399 15306
rect 7451 15254 7610 15306
rect 7662 15254 7738 15306
rect 6451 14843 7738 15254
rect 6451 14791 6766 14843
rect 6818 14791 6977 14843
rect 7029 14791 7188 14843
rect 7240 14791 7399 14843
rect 7451 14791 7610 14843
rect 7662 14791 7738 14843
rect 6451 14413 7738 14791
rect 8186 14845 9066 14884
rect 8186 14789 8222 14845
rect 8278 14789 8433 14845
rect 8489 14789 8644 14845
rect 8700 14789 8855 14845
rect 8911 14789 9066 14845
rect 8186 14413 9066 14789
rect 9591 14413 10186 15401
rect 10276 15074 10941 15401
rect 10276 15022 10376 15074
rect 10428 15022 10587 15074
rect 10639 15022 10798 15074
rect 10850 15022 10941 15074
rect 10276 14413 10941 15022
rect 11537 15331 11846 15401
rect 13994 15378 14545 15419
rect 11537 15328 11575 15331
rect 11627 15328 11755 15331
rect 11807 15328 11846 15331
rect 11537 15272 11573 15328
rect 11629 15272 11753 15328
rect 11809 15272 11846 15328
rect 11537 15113 11846 15272
rect 13531 15317 13871 15358
rect 13531 15265 13569 15317
rect 13621 15265 13781 15317
rect 13833 15265 13871 15317
rect 13531 15224 13871 15265
rect 13994 15326 14033 15378
rect 14085 15326 14244 15378
rect 14296 15326 14455 15378
rect 14507 15326 14545 15378
rect 11537 15061 11575 15113
rect 11627 15061 11755 15113
rect 11807 15061 11846 15113
rect 11537 14413 11846 15061
rect 12294 14845 13478 14884
rect 12294 14789 12331 14845
rect 12387 14789 12542 14845
rect 12598 14789 12753 14845
rect 12809 14789 12964 14845
rect 13020 14789 13175 14845
rect 13231 14789 13385 14845
rect 13441 14789 13478 14845
rect 12294 14750 13478 14789
rect 13994 14838 14545 15326
rect 13994 14782 14031 14838
rect 14087 14782 14242 14838
rect 14298 14782 14453 14838
rect 14509 14782 14545 14838
rect 13994 14744 14545 14782
rect 15026 15378 15887 15419
rect 15026 15326 15100 15378
rect 15152 15326 15311 15378
rect 15363 15326 15522 15378
rect 15574 15326 15733 15378
rect 15785 15326 15887 15378
rect 12040 14428 12639 14564
rect 12040 14372 12100 14428
rect 12156 14372 12311 14428
rect 12367 14372 12522 14428
rect 12578 14372 12639 14428
rect 15026 14413 15887 15326
rect 20112 15306 21313 15401
rect 20112 15254 20151 15306
rect 20203 15254 20362 15306
rect 20414 15254 20573 15306
rect 20625 15254 20784 15306
rect 20836 15254 21313 15306
rect 20112 14843 21313 15254
rect 20112 14791 20151 14843
rect 20203 14791 20362 14843
rect 20414 14791 20573 14843
rect 20625 14791 20784 14843
rect 20836 14791 21313 14843
rect 20112 14413 21313 14791
rect 21421 15328 22236 15419
rect 21421 15272 21458 15328
rect 21514 15272 21669 15328
rect 21725 15272 21880 15328
rect 21936 15272 22091 15328
rect 22147 15272 22236 15328
rect 21421 14413 22236 15272
rect 22365 14845 23338 14884
rect 22365 14789 22402 14845
rect 22458 14789 22613 14845
rect 22669 14789 22824 14845
rect 22880 14789 23035 14845
rect 23091 14789 23246 14845
rect 23302 14789 23338 14845
rect 22365 14751 23338 14789
rect 23549 14413 25677 15476
rect 12040 14299 12639 14372
rect 8561 -21 8691 112
rect 12841 -164 12971 -31
rect 13219 -164 13348 -31
rect 13597 -164 13726 -31
rect 13974 -164 14104 -31
rect 14352 -164 14481 -31
rect 14730 -164 14859 -31
rect 16882 -164 17011 -31
rect 17260 -164 17389 -31
rect 17637 -164 17767 -31
rect 18015 -164 18144 -31
rect 18393 -164 18522 -31
rect 18770 -164 18900 -31
rect 19148 -164 19277 -31
rect 19526 -164 19655 -31
<< via2 >>
rect 5611 15272 5667 15328
rect 5822 15272 5878 15328
rect 6033 15272 6089 15328
rect 6244 15272 6300 15328
rect 4371 14845 4427 14847
rect 4371 14793 4373 14845
rect 4373 14793 4425 14845
rect 4425 14793 4427 14845
rect 4371 14791 4427 14793
rect 4582 14845 4638 14847
rect 4582 14793 4584 14845
rect 4584 14793 4636 14845
rect 4636 14793 4638 14845
rect 4582 14791 4638 14793
rect 4793 14845 4849 14847
rect 4793 14793 4795 14845
rect 4795 14793 4847 14845
rect 4847 14793 4849 14845
rect 4793 14791 4849 14793
rect 5004 14845 5060 14847
rect 5004 14793 5006 14845
rect 5006 14793 5058 14845
rect 5058 14793 5060 14845
rect 5004 14791 5060 14793
rect 5215 14845 5271 14847
rect 5215 14793 5217 14845
rect 5217 14793 5269 14845
rect 5269 14793 5271 14845
rect 5215 14791 5271 14793
rect 8222 14789 8278 14845
rect 8433 14789 8489 14845
rect 8644 14789 8700 14845
rect 8855 14789 8911 14845
rect 11573 15279 11575 15328
rect 11575 15279 11627 15328
rect 11627 15279 11629 15328
rect 11573 15272 11629 15279
rect 11753 15279 11755 15328
rect 11755 15279 11807 15328
rect 11807 15279 11809 15328
rect 11753 15272 11809 15279
rect 12331 14843 12387 14845
rect 12331 14791 12333 14843
rect 12333 14791 12385 14843
rect 12385 14791 12387 14843
rect 12331 14789 12387 14791
rect 12542 14843 12598 14845
rect 12542 14791 12544 14843
rect 12544 14791 12596 14843
rect 12596 14791 12598 14843
rect 12542 14789 12598 14791
rect 12753 14843 12809 14845
rect 12753 14791 12755 14843
rect 12755 14791 12807 14843
rect 12807 14791 12809 14843
rect 12753 14789 12809 14791
rect 12964 14843 13020 14845
rect 12964 14791 12966 14843
rect 12966 14791 13018 14843
rect 13018 14791 13020 14843
rect 12964 14789 13020 14791
rect 13175 14843 13231 14845
rect 13175 14791 13177 14843
rect 13177 14791 13229 14843
rect 13229 14791 13231 14843
rect 13175 14789 13231 14791
rect 13385 14843 13441 14845
rect 13385 14791 13387 14843
rect 13387 14791 13439 14843
rect 13439 14791 13441 14843
rect 13385 14789 13441 14791
rect 14031 14782 14087 14838
rect 14242 14782 14298 14838
rect 14453 14782 14509 14838
rect 12100 14372 12156 14428
rect 12311 14372 12367 14428
rect 12522 14372 12578 14428
rect 21458 15272 21514 15328
rect 21669 15272 21725 15328
rect 21880 15272 21936 15328
rect 22091 15272 22147 15328
rect 22402 14843 22458 14845
rect 22402 14791 22404 14843
rect 22404 14791 22456 14843
rect 22456 14791 22458 14843
rect 22402 14789 22458 14791
rect 22613 14843 22669 14845
rect 22613 14791 22615 14843
rect 22615 14791 22667 14843
rect 22667 14791 22669 14843
rect 22613 14789 22669 14791
rect 22824 14843 22880 14845
rect 22824 14791 22826 14843
rect 22826 14791 22878 14843
rect 22878 14791 22880 14843
rect 22824 14789 22880 14791
rect 23035 14843 23091 14845
rect 23035 14791 23037 14843
rect 23037 14791 23089 14843
rect 23089 14791 23091 14843
rect 23035 14789 23091 14791
rect 23246 14843 23302 14845
rect 23246 14791 23248 14843
rect 23248 14791 23300 14843
rect 23300 14791 23302 14843
rect 23246 14789 23302 14791
<< metal3 >>
rect 69 15233 199 15367
rect 1725 15328 25945 15401
rect 1725 15272 5611 15328
rect 5667 15272 5822 15328
rect 5878 15272 6033 15328
rect 6089 15272 6244 15328
rect 6300 15272 11573 15328
rect 11629 15272 11753 15328
rect 11809 15272 21458 15328
rect 21514 15272 21669 15328
rect 21725 15272 21880 15328
rect 21936 15272 22091 15328
rect 22147 15272 25945 15328
rect 1725 15199 25945 15272
rect -1 14773 128 14907
rect 1725 14847 5307 14941
rect 1725 14791 4371 14847
rect 4427 14791 4582 14847
rect 4638 14791 4793 14847
rect 4849 14791 5004 14847
rect 5060 14791 5215 14847
rect 5271 14791 5307 14847
rect 1725 14739 5307 14791
rect 8186 14845 13478 14884
rect 8186 14789 8222 14845
rect 8278 14789 8433 14845
rect 8489 14789 8644 14845
rect 8700 14789 8855 14845
rect 8911 14789 12331 14845
rect 12387 14789 12542 14845
rect 12598 14789 12753 14845
rect 12809 14789 12964 14845
rect 13020 14789 13175 14845
rect 13231 14789 13385 14845
rect 13441 14789 13478 14845
rect 13994 14838 14545 14877
rect 13994 14803 14031 14838
rect 8186 14750 13478 14789
rect 13993 14782 14031 14803
rect 14087 14782 14242 14838
rect 14298 14782 14453 14838
rect 14509 14782 14545 14838
rect 13993 14744 14545 14782
rect 22365 14845 25945 14941
rect 22365 14789 22402 14845
rect 22458 14789 22613 14845
rect 22669 14789 22824 14845
rect 22880 14789 23035 14845
rect 23091 14789 23246 14845
rect 23302 14789 25945 14845
rect 69 14333 199 14467
rect 12063 14428 12615 14467
rect 13993 14432 14092 14744
rect 22365 14739 25945 14789
rect 27640 14773 27769 14907
rect 12063 14372 12100 14428
rect 12156 14372 12311 14428
rect 12367 14372 12522 14428
rect 12578 14372 12615 14428
rect 12063 14333 12615 14372
rect -1 13873 128 14027
rect 27640 13873 27769 14007
rect -1 12993 128 13127
rect 27640 12993 27769 13127
rect -1 12073 128 12207
rect 27640 12073 27769 12207
rect -1 11193 128 11327
rect 27640 11193 27769 11327
rect -1 10273 128 10407
rect 27640 10273 27769 10407
rect -1 9393 128 9527
rect 27640 9393 27769 9527
rect -1 8473 128 8607
rect 27640 8473 27769 8607
rect -1 7593 128 7727
rect 27640 7593 27769 7727
rect -1 6673 128 6807
rect 27640 6673 27769 6807
rect -1 5793 128 5927
rect 27640 5793 27769 5927
rect -1 4873 128 5007
rect 27640 4873 27769 5007
rect -1 3993 128 4127
rect 27640 3993 27769 4127
rect -1 3073 128 3207
rect 27640 3073 27769 3207
rect -1 2193 128 2327
rect 27640 2193 27769 2327
rect -1 1273 128 1407
rect 27640 1273 27769 1407
rect -1 393 128 527
rect 27640 393 27769 527
use M1_NACTIVE$$203393068_128x8m81  M1_NACTIVE$$203393068_128x8m81_0
timestamp 1666464484
transform 1 0 14063 0 1 15359
box 0 0 1 1
use M1_NWELL$$204218412_128x8m81  M1_NWELL$$204218412_128x8m81_0
timestamp 1666464484
transform -1 0 25568 0 1 15286
box -221 -717 1960 228
use M1_NWELL$$204218412_128x8m81  M1_NWELL$$204218412_128x8m81_1
timestamp 1666464484
transform 1 0 2200 0 1 15286
box -221 -717 1960 228
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_0
timestamp 1666464484
transform 1 0 11463 0 1 15359
box -78 -80 1817 80
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_1
timestamp 1666464484
transform 1 0 21475 0 1 15359
box -78 -80 1817 80
use M1_PACTIVE$$204148780_128x8m81  M1_PACTIVE$$204148780_128x8m81_2
timestamp 1666464484
transform 1 0 4390 0 1 15359
box -78 -80 1817 80
use M1_PACTIVE$$204149804_128x8m81  M1_PACTIVE$$204149804_128x8m81_0
timestamp 1666464484
transform 1 0 15860 0 1 15359
box 0 0 1 1
use M1_POLY2$$204150828_128x8m81  M1_POLY2$$204150828_128x8m81_0
timestamp 1666464484
transform 1 0 9381 0 1 15048
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1666464484
transform 1 0 15413 0 1 15341
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_0
timestamp 1666464484
transform 0 -1 13712 1 0 15293
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_1
timestamp 1666464484
transform 1 0 15625 0 1 15001
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_2
timestamp 1666464484
transform 1 0 18313 0 1 15036
box 0 0 1 1
use M1_POLY24310590548739_128x8m81  M1_POLY24310590548739_128x8m81_3
timestamp 1666464484
transform 1 0 12040 0 1 14961
box 0 0 1 1
use M2_M1$$201262124_128x8m81  M2_M1$$201262124_128x8m81_0
timestamp 1666464484
transform 1 0 13701 0 1 15291
box 0 0 1 1
use M2_M1$$204138540_128x8m81  M2_M1$$204138540_128x8m81_0
timestamp 1666464484
transform 1 0 10402 0 1 15048
box 0 0 1 1
use M2_M1$$204138540_128x8m81  M2_M1$$204138540_128x8m81_1
timestamp 1666464484
transform 1 0 14059 0 1 15352
box 0 0 1 1
use M2_M1$$204139564_128x8m81  M2_M1$$204139564_128x8m81_0
timestamp 1666464484
transform 1 0 11601 0 1 15305
box 0 0 1 1
use M2_M1$$204140588_128x8m81  M2_M1$$204140588_128x8m81_0
timestamp 1666464484
transform 1 0 12359 0 1 14817
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_0
timestamp 1666464484
transform 1 0 15126 0 1 15352
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_1
timestamp 1666464484
transform 1 0 20177 0 1 15280
box 0 0 1 1
use M2_M1$$204141612_128x8m81  M2_M1$$204141612_128x8m81_2
timestamp 1666464484
transform 1 0 20177 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_0
timestamp 1666464484
transform 1 0 6792 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_1
timestamp 1666464484
transform 1 0 22430 0 1 14817
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_2
timestamp 1666464484
transform 1 0 4399 0 1 14819
box 0 0 1 1
use M2_M1$$204220460_128x8m81  M2_M1$$204220460_128x8m81_3
timestamp 1666464484
transform 1 0 6792 0 1 15280
box 0 0 1 1
use M2_M1$$204221484_128x8m81  M2_M1$$204221484_128x8m81_0
timestamp 1666464484
transform -1 0 25612 0 1 15300
box -65 -502 1751 67
use M2_M1$$204221484_128x8m81  M2_M1$$204221484_128x8m81_1
timestamp 1666464484
transform 1 0 2156 0 1 15300
box -65 -502 1751 67
use M2_M1$$204222508_128x8m81  M2_M1$$204222508_128x8m81_0
timestamp 1666464484
transform 1 0 21486 0 1 15300
box -65 -284 697 67
use M2_M1$$204222508_128x8m81  M2_M1$$204222508_128x8m81_1
timestamp 1666464484
transform 1 0 5639 0 1 15300
box -65 -284 697 67
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_0
timestamp 1666464484
transform 1 0 5639 0 1 15300
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_1
timestamp 1666464484
transform 1 0 8250 0 1 14817
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_2
timestamp 1666464484
transform 1 0 21486 0 1 15300
box 0 0 1 1
use M3_M2$$204142636_128x8m81  M3_M2$$204142636_128x8m81_3
timestamp 1666464484
transform 1 0 21486 0 1 15300
box 0 0 1 1
use M3_M2$$204143660_128x8m81  M3_M2$$204143660_128x8m81_0
timestamp 1666464484
transform 1 0 11601 0 1 15300
box 0 0 1 1
use M3_M2$$204144684_128x8m81  M3_M2$$204144684_128x8m81_0
timestamp 1666464484
transform 1 0 22430 0 1 14817
box 0 0 1 1
use M3_M2$$204144684_128x8m81  M3_M2$$204144684_128x8m81_1
timestamp 1666464484
transform 1 0 4399 0 1 14819
box 0 0 1 1
use M3_M2$$204145708_128x8m81  M3_M2$$204145708_128x8m81_0
timestamp 1666464484
transform 1 0 12359 0 1 14817
box 0 0 1 1
use M3_M2$$204146732_128x8m81  M3_M2$$204146732_128x8m81_0
timestamp 1666464484
transform 1 0 14059 0 1 14810
box 0 0 1 1
use M3_M2$$204147756_128x8m81  M3_M2$$204147756_128x8m81_0
timestamp 1666464484
transform 1 0 12339 0 1 14400
box 0 0 1 1
use nmos_1p2$$204213292_R90_128x8m81  nmos_1p2$$204213292_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 6346 1 0 14903
box -119 -71 177 2091
use nmos_1p2$$204215340_128x8m81  nmos_1p2$$204215340_128x8m81_0
timestamp 1666464484
transform 0 -1 13604 -1 0 14962
box -119 -71 177 1389
use nmos_5p04310590548799_128x8m81  nmos_5p04310590548799_128x8m81_0
timestamp 1666464484
transform 0 -1 23346 1 0 14872
box -88 -44 208 2066
use nmos_5p043105905487111_128x8m81  nmos_5p043105905487111_128x8m81_0
timestamp 1666464484
transform 0 -1 16283 1 0 14872
box -88 -44 208 572
use nmos_5p043105905487111_128x8m81  nmos_5p043105905487111_128x8m81_1
timestamp 1666464484
transform 0 -1 11913 1 0 14872
box -88 -44 208 572
use pmos_1p2$$204216364_128x8m81  pmos_1p2$$204216364_128x8m81_0
timestamp 1666464484
transform 0 -1 20950 1 0 14903
box -296 -137 586 2646
use pmos_1p2$$204216364_128x8m81  pmos_1p2$$204216364_128x8m81_1
timestamp 1666464484
transform 0 -1 9245 1 0 14903
box -296 -137 586 2646
use pmos_1p2$$204217388_R90_128x8m81  pmos_1p2$$204217388_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 11004 1 0 14903
box -295 -137 355 1454
use pmos_5p043105905487100_128x8m81  pmos_5p043105905487100_128x8m81_0
timestamp 1666464484
transform 0 -1 15304 1 0 14872
box -208 -120 328 1438
use pmos_5p043105905487100_128x8m81  pmos_5p043105905487100_128x8m81_1
timestamp 1666464484
transform 0 -1 17974 1 0 14872
box -208 -120 328 1438
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_0
timestamp 1666464484
transform 0 -1 2203 -1 0 14550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_1
timestamp 1666464484
transform 0 -1 2203 -1 0 12750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_2
timestamp 1666464484
transform 0 -1 2203 -1 0 10950
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_3
timestamp 1666464484
transform 0 -1 2203 -1 0 9150
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_4
timestamp 1666464484
transform 0 -1 2203 -1 0 7350
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_5
timestamp 1666464484
transform 0 -1 2203 -1 0 5550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_6
timestamp 1666464484
transform 0 -1 2203 -1 0 3750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_7
timestamp 1666464484
transform 0 -1 2203 -1 0 1950
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_8
timestamp 1666464484
transform 0 1 25566 -1 0 14550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_9
timestamp 1666464484
transform 0 1 25566 -1 0 12750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_10
timestamp 1666464484
transform 0 1 25566 -1 0 10950
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_11
timestamp 1666464484
transform 0 1 25566 -1 0 9150
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_12
timestamp 1666464484
transform 0 1 25566 -1 0 7350
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_13
timestamp 1666464484
transform 0 1 25566 -1 0 5550
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_14
timestamp 1666464484
transform 0 1 25566 -1 0 3750
box -60 -407 2159 5567
use pmoscap_W2_5_477_R270_128x8m81  pmoscap_W2_5_477_R270_128x8m81_15
timestamp 1666464484
transform 0 1 25566 -1 0 1950
box -60 -407 2159 5567
use pmoscap_W2_5_R270_128x8m81  pmoscap_W2_5_R270_128x8m81_0
timestamp 1666464484
transform 0 -1 2203 -1 0 15450
box -60 -407 1259 3251
use pmoscap_W2_5_R270_128x8m81  pmoscap_W2_5_R270_128x8m81_1
timestamp 1666464484
transform 0 1 25566 -1 0 15450
box -60 -407 1259 3251
use xdec16_128x8_128x8m81  xdec16_128x8_128x8m81_0
timestamp 1666464484
transform 1 0 1726 0 1 0
box 0 -228 24219 14628
<< labels >>
rlabel metal3 s 27705 14840 27705 14840 4 DRWL
port 1 nsew
rlabel metal3 s 27705 5860 27705 5860 4 RWL[6]
port 2 nsew
rlabel metal3 s 27705 4060 27705 4060 4 RWL[4]
port 3 nsew
rlabel metal3 s 27705 2260 27705 2260 4 RWL[2]
port 4 nsew
rlabel metal3 s 27705 460 27705 460 4 RWL[0]
port 5 nsew
rlabel metal3 s 27705 1340 27705 1340 4 RWL[1]
port 6 nsew
rlabel metal3 s 27705 3140 27705 3140 4 RWL[3]
port 7 nsew
rlabel metal3 s 27705 4940 27705 4940 4 RWL[5]
port 8 nsew
rlabel metal3 s 27705 6740 27705 6740 4 RWL[7]
port 9 nsew
rlabel metal3 s 27705 7660 27705 7660 4 RWL[8]
port 10 nsew
rlabel metal3 s 27705 8540 27705 8540 4 RWL[9]
port 11 nsew
rlabel metal3 s 27705 9460 27705 9460 4 RWL[10]
port 12 nsew
rlabel metal3 s 27705 10340 27705 10340 4 RWL[11]
port 13 nsew
rlabel metal3 s 27705 11260 27705 11260 4 RWL[12]
port 14 nsew
rlabel metal3 s 27705 12140 27705 12140 4 RWL[13]
port 15 nsew
rlabel metal3 s 27705 13060 27705 13060 4 RWL[14]
port 16 nsew
rlabel metal3 s 27705 13940 27705 13940 4 RWL[15]
port 17 nsew
rlabel metal3 s 64 9460 64 9460 4 LWL[10]
port 18 nsew
rlabel metal3 s 64 10340 64 10340 4 LWL[11]
port 19 nsew
rlabel metal3 s 64 11260 64 11260 4 LWL[12]
port 20 nsew
rlabel metal3 s 64 12140 64 12140 4 LWL[13]
port 21 nsew
rlabel metal3 s 64 13060 64 13060 4 LWL[14]
port 22 nsew
rlabel metal3 s 64 13940 64 13940 4 LWL[15]
port 23 nsew
rlabel metal3 s 64 4940 64 4940 4 LWL[5]
port 24 nsew
rlabel metal3 s 64 4060 64 4060 4 LWL[4]
port 25 nsew
rlabel metal3 s 64 3140 64 3140 4 LWL[3]
port 26 nsew
rlabel metal3 s 64 2260 64 2260 4 LWL[2]
port 27 nsew
rlabel metal3 s 64 1340 64 1340 4 LWL[1]
port 28 nsew
rlabel metal3 s 64 460 64 460 4 LWL[0]
port 29 nsew
rlabel metal3 s 64 7660 64 7660 4 LWL[8]
port 30 nsew
rlabel metal3 s 64 8540 64 8540 4 LWL[9]
port 31 nsew
rlabel metal3 s 64 5860 64 5860 4 LWL[6]
port 32 nsew
rlabel metal3 s 64 6740 64 6740 4 LWL[7]
port 33 nsew
rlabel metal3 s 134 15300 134 15300 4 vss
port 34 nsew
rlabel metal3 s 134 14400 134 14400 4 vdd
port 35 nsew
rlabel metal3 s 64 14840 64 14840 4 DLWL
port 36 nsew
rlabel metal2 s 14794 -97 14794 -97 4 xb[0]
port 37 nsew
rlabel metal2 s 14417 -97 14417 -97 4 xb[1]
port 38 nsew
rlabel metal2 s 14039 -97 14039 -97 4 xb[2]
port 39 nsew
rlabel metal2 s 13661 -97 13661 -97 4 xb[3]
port 40 nsew
rlabel metal2 s 16947 -97 16947 -97 4 xa[7]
port 41 nsew
rlabel metal2 s 17324 -97 17324 -97 4 xa[6]
port 42 nsew
rlabel metal2 s 17702 -97 17702 -97 4 xa[5]
port 43 nsew
rlabel metal2 s 18080 -97 18080 -97 4 xa[4]
port 44 nsew
rlabel metal2 s 19591 -97 19591 -97 4 xa[0]
port 45 nsew
rlabel metal2 s 8626 45 8626 45 4 men
port 46 nsew
rlabel metal2 s 18457 -97 18457 -97 4 xa[3]
port 47 nsew
rlabel metal2 s 18835 -97 18835 -97 4 xa[2]
port 48 nsew
rlabel metal2 s 19213 -97 19213 -97 4 xa[1]
port 49 nsew
rlabel metal2 s 13284 -97 13284 -97 4 xc[0]
port 50 nsew
rlabel metal2 s 12906 -97 12906 -97 4 xc[1]
port 51 nsew
<< properties >>
string GDS_END 2206640
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 2192530
<< end >>
