magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 448 844
rect 69 469 115 724
rect 49 60 95 232
rect 244 106 319 330
rect 0 -60 448 60
<< obsm1 >>
rect 273 437 319 678
rect 174 390 319 437
<< labels >>
rlabel metal1 s 244 106 319 330 6 ZN
port 1 nsew default output
rlabel metal1 s 0 724 448 844 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 69 469 115 724 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 49 60 95 232 6 VSS
port 3 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 448 60 8 VSS
port 3 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 448 784
string LEFclass core TIELOW
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 314166
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 312208
<< end >>
