* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addf_1 A B CI CO S VDD VSS
X0 a_1072_215# a_952_171# a_124_53# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 VSS B a_1904_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 VSS CI a_1072_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 VDD B a_1924_573# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X4 VSS a_124_53# S & Metric 1.00 nmos_6p0 w=1.18u l=0.6u
X5 a_124_53# CI a_680_594# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X6 VDD A a_2764_573# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X7 a_952_171# CI a_1904_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_1924_573# A VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X9 CO a_952_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_680_594# B a_512_594# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X11 a_2764_573# B a_952_171# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X12 a_124_53# CI a_680_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 VDD A a_1072_594# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X14 CO a_952_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_1072_215# B VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 VDD a_124_53# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_680_215# B a_512_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 a_1904_215# A VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 VSS A a_2784_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X20 VSS A a_1072_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 a_512_215# A VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_1072_594# a_952_171# a_124_53# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X23 a_512_594# A VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X24 a_1072_594# B VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X25 a_952_171# CI a_1924_573# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X26 a_2784_215# B a_952_171# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 VDD CI a_1072_594# w_n86_453# pmos_6p0 w=0.99u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addf_2 A B CI CO S VDD VSS
X0 VDD A a_3016_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X1 S a_132_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD a_132_25# S w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VDD A a_1284_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X4 a_1184_129# CI a_2136_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X5 VSS a_1184_129# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1284_573# B VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X7 VDD CI a_1284_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X8 a_3016_573# B a_1184_129# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X9 a_132_25# CI a_912_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 VSS A a_3016_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X11 a_2136_573# A VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X12 a_1184_129# CI a_2136_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X13 a_1304_173# B VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X14 a_912_173# B a_744_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X15 a_132_25# CI a_912_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X16 a_2136_173# A VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 a_764_573# A VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X18 CO a_1184_129# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 VDD B a_2136_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X20 a_3016_173# B a_1184_129# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X21 S a_132_25# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X22 a_1284_573# a_1184_129# a_132_25# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X23 VSS a_132_25# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 VDD a_1184_129# CO w_n86_453# pmos_6p0 w=1.8u l=0.5u
X25 VSS A a_1304_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X26 CO a_1184_129# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_744_173# A VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X28 a_1304_173# a_1184_129# a_132_25# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X29 VSS B a_2136_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X30 VSS CI a_1304_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X31 a_912_573# B a_764_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addf_4 A B CI CO S VDD VSS
X0 a_1760_573# a_1640_129# a_140_25# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X1 VDD B a_2612_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X2 a_1200_573# A VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X3 a_3452_573# B a_1640_129# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X4 VSS A a_3472_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X5 CO a_1640_129# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_2612_573# A VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X7 CO a_1640_129# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_140_25# CI a_1368_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X9 a_3472_173# B a_1640_129# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 S a_140_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 S a_140_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VDD CI a_1760_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X13 CO a_1640_129# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_2592_173# A VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X15 VSS a_1640_129# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1368_173# B a_1200_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 VSS A a_1760_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X18 VSS a_1640_129# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VDD a_140_25# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 a_140_25# CI a_1368_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X21 a_1760_573# B VDD w_n86_453# pmos_6p0 w=1.39u l=0.5u
X22 a_1640_129# CI a_2612_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X23 VSS B a_2592_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X24 a_1200_173# A VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X25 VSS CI a_1760_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X26 VDD a_140_25# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 a_1368_573# B a_1200_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X28 VDD A a_1760_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X29 S a_140_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_1760_173# B VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X31 a_1640_129# CI a_2592_173# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X32 VDD a_1640_129# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 a_1760_173# a_1640_129# a_140_25# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X34 VDD A a_3452_573# w_n86_453# pmos_6p0 w=1.39u l=0.5u
X35 VDD a_1640_129# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 VSS a_140_25# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 CO a_1640_129# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 S a_140_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 VSS a_140_25# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addf_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addh_1 A B CO S VDD VSS
X0 a_1052_691# B VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 a_844_201# A a_1052_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 a_1052_201# A a_1052_691# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_124_25# B a_516_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 S a_1052_201# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_516_201# A VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 a_124_25# A VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X7 a_1052_201# B a_844_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X8 VDD a_124_25# a_1052_201# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X9 S a_1052_201# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD a_124_25# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS a_124_25# a_844_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X12 VSS a_124_25# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD B a_124_25# w_n86_453# pmos_6p0 w=0.915u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addh_2 A B CO S VDD VSS
X0 a_128_25# A VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_1248_69# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD B a_128_25# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_128_25# B a_696_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD a_128_25# a_1248_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD a_128_25# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_1040_69# A a_1248_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_1248_69# A a_1248_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD a_1248_69# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_1248_573# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 S a_1248_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_696_69# A VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 CO a_128_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 CO a_128_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 S a_1248_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VSS a_128_25# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VSS a_128_25# a_1040_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_1248_69# B a_1040_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__addh_4 A B CO S VDD VSS
X0 VDD B a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_1106_573# A a_1778_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A a_672_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD a_234_573# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_672_68# B a_234_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_1106_573# A a_1116_156# & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X6 a_1116_156# a_234_573# VSS & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X7 a_1778_573# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_1320_573# A a_1106_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 CO a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD a_234_573# CO w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_1106_573# B a_1116_156# & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X12 VDD a_234_573# a_1106_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_1106_573# a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VDD a_1106_573# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_244_68# A VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VSS a_234_573# a_1116_156# & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X17 VSS a_1106_573# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD B a_1320_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS a_1106_573# S & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 CO a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_1116_156# B a_1106_573# & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X22 VSS a_234_573# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 CO a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_234_573# B a_244_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 CO a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 S a_1106_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_234_573# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 S a_1106_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 VDD a_1106_573# S w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 a_1116_156# A a_1106_573# & Metric 1.00 nmos_6p0 w=0.88u l=0.6u
X31 S a_1106_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 S a_1106_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 a_234_573# A VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 VDD A a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VSS a_234_573# CO & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__addh_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1 A1 A2 VDD VSS Z
X0 Z a_36_201# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS A2 a_244_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 a_36_201# A1 VDD w_n86_453# pmos_6p0 w=0.82u l=0.5u
X3 VDD A2 a_36_201# w_n86_453# pmos_6p0 w=0.82u l=0.5u
X4 a_244_201# A1 a_36_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 Z a_36_201# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_2 A1 A2 VDD VSS Z
X0 VSS A2 a_247_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 Z a_39_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS a_39_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD a_39_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_247_69# A1 a_39_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_39_69# A1 VDD w_n86_453# pmos_6p0 w=1.64u l=0.5u
X6 VDD A2 a_39_69# w_n86_453# pmos_6p0 w=1.64u l=0.5u
X7 Z a_39_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_4 A1 A2 VDD VSS Z
X0 a_224_611# A2 VDD w_n86_453# pmos_6p0 w=1.64u l=0.5u
X1 VDD a_224_611# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A2 a_659_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 Z a_224_611# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VDD A1 a_224_611# w_n86_453# pmos_6p0 w=1.64u l=0.5u
X5 a_224_611# A1 VDD w_n86_453# pmos_6p0 w=1.64u l=0.5u
X6 VDD a_224_611# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 Z a_224_611# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD A2 a_224_611# w_n86_453# pmos_6p0 w=1.64u l=0.5u
X9 Z a_224_611# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VSS a_224_611# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_224_611# A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_659_69# A1 a_224_611# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VSS a_224_611# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 Z a_224_611# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and3_1 A1 A2 A3 VDD VSS Z
X0 a_36_201# A2 VDD w_n86_453# pmos_6p0 w=0.73u l=0.5u
X1 VDD A3 a_36_201# w_n86_453# pmos_6p0 w=0.73u l=0.5u
X2 a_428_201# A2 a_244_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X3 VSS A3 a_428_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_244_201# A1 a_36_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 Z a_36_201# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 Z a_36_201# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD A1 a_36_201# w_n86_453# pmos_6p0 w=0.73u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and3_2 A1 A2 A3 VDD VSS Z
X0 VDD A1 a_47_69# w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 a_47_69# A2 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 VDD A3 a_47_69# w_n86_453# pmos_6p0 w=1.46u l=0.5u
X3 Z a_47_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_47_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS a_47_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD a_47_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS A3 a_439_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_255_69# A1 a_47_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_439_69# A2 a_255_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and3_4 A1 A2 A3 VDD VSS Z
X0 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_224_573# A3 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD A2 a_224_573# w_n86_453# pmos_6p0 w=1.46u l=0.5u
X4 a_260_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS A3 a_1040_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_224_573# A1 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X7 a_856_69# A1 a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD A1 a_224_573# w_n86_453# pmos_6p0 w=1.46u l=0.5u
X10 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_224_573# A2 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X13 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_224_573# A1 a_428_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD A3 a_224_573# w_n86_453# pmos_6p0 w=1.46u l=0.5u
X16 a_428_69# A2 a_260_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_1040_69# A2 a_856_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and3_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and4_1 A1 A2 A3 A4 VDD VSS Z
X0 a_440_201# A2 a_256_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 a_48_201# A1 VDD w_n86_453# pmos_6p0 w=0.64u l=0.5u
X2 VDD A2 a_48_201# w_n86_453# pmos_6p0 w=0.64u l=0.5u
X3 a_644_201# A3 a_440_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_48_201# A3 VDD w_n86_453# pmos_6p0 w=0.64u l=0.5u
X5 VSS A4 a_644_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 VDD A4 a_48_201# w_n86_453# pmos_6p0 w=0.64u l=0.5u
X7 a_256_201# A1 a_48_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X8 Z a_48_201# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 Z a_48_201# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and4_2 A1 A2 A3 A4 VDD VSS Z
X0 VSS A4 a_643_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 Z a_47_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_47_69# A1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X3 VDD A2 a_47_69# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X4 a_47_69# A3 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X5 VDD A4 a_47_69# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X6 Z a_47_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_643_69# A3 a_439_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD a_47_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_255_69# A1 a_47_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_439_69# A2 a_255_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS a_47_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__and4_4 A1 A2 A3 A4 VDD VSS Z
X0 VDD A1 a_227_573# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X1 a_1247_69# A2 a_1063_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 Z a_227_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_227_573# A1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X4 Z a_227_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_1063_69# A1 a_227_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD a_227_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS a_227_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_431_69# A3 a_247_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS A4 a_1451_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VDD A2 a_227_573# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X11 a_227_573# A3 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X12 VSS a_227_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD A4 a_227_573# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X14 a_635_69# A2 a_431_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_247_69# A4 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_227_573# A4 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X17 VDD A3 a_227_573# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X18 Z a_227_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_227_573# A2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X20 a_227_573# A1 a_635_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 a_1451_69# A3 a_1247_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD a_227_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 Z a_227_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__and4_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__antenna.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__antenna I VDD VSS
D0 & Metric 1.00 I np_6p0 pj=1.85u area=0.2034p
D1 I w_n86_453# pn_6p0 pj=1.85u area=0.2034p
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__antenna.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_1 A1 A2 B VDD VSS ZN
X0 ZN A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD B a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 ZN A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS B ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_2 A1 A2 B VDD VSS ZN
X0 a_49_573# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN A2 a_49_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS B ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X3 ZN A1 a_741_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_1133_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS A2 a_1133_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_49_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VDD B a_49_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A1 a_49_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_741_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN B VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X11 a_49_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi21_4 A1 A2 B VDD VSS ZN
X0 a_288_68# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_1072_68# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_76_574# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 ZN A1 a_288_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN A1 a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_76_574# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_76_574# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_680_68# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS B ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X9 VDD B a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD B a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_76_574# B VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS B ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X13 ZN A2 a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_76_574# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_1464_68# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 ZN B VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X17 ZN A1 a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VSS A2 a_1464_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS A2 a_680_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_76_574# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 ZN B VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X22 ZN A2 a_76_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 ZN A1 a_1072_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi21_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_1 A1 A2 B1 B2 VDD VSS ZN
X0 a_665_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS A2 a_665_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN B1 a_257_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD B2 a_49_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_49_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A1 a_49_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_49_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_257_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_2 A1 A2 B1 B2 VDD VSS ZN
X0 VSS B2 a_659_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN A1 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD B2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_1060_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_36_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD B1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS A2 a_1468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_36_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_659_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_1468_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 ZN A1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_36_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi22_4 A1 A2 B1 B2 VDD VSS ZN
X0 a_652_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS B2 a_652_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A1 a_1924_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN B1 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD B2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS A2 a_3148_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1060_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_36_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD B1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS B2 a_1468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_2332_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_36_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS A2 a_2332_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD B2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN A1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_3148_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 ZN A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN A1 a_2740_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_2740_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_36_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_36_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 ZN A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 ZN A1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 a_1468_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 VDD B1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_36_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_36_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_1924_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi22_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_1 A1 A2 B C VDD VSS ZN
X0 a_653_573# B a_37_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 ZN A2 a_37_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS B ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 a_37_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD C a_653_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_245_96# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X7 ZN A1 a_245_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_2 A1 A2 B C VDD VSS ZN
X0 a_636_70# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X1 ZN A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A2 a_636_70# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X3 a_36_573# B a_1492_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS B ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 ZN A1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_244_70# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X9 a_36_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN A1 a_244_70# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X11 a_1492_573# C VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1124_573# B a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 VDD C a_1124_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN B VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi211_4 A1 A2 B C VDD VSS ZN
X0 ZN A1 a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_3638_573# C VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN B VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 a_170_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_786_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X6 ZN A2 a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1194_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X8 ZN A1 a_1194_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X9 VDD C a_2042_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_170_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X12 ZN A1 a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_170_573# B a_2574_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN A1 a_368_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X15 VSS A2 a_1602_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X16 VSS B ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X17 VDD C a_3106_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_1602_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X19 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_170_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_170_573# B a_3638_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 VSS B ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 VSS A2 a_786_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X24 a_368_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X25 ZN A2 a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_2574_573# C VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 a_170_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X29 a_3106_573# B a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 a_2042_573# B a_170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 ZN B VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi211_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_1 A1 A2 B1 B2 C VDD VSS ZN
X0 a_252_96# B2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X1 ZN B1 a_252_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X2 a_940_96# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X3 a_660_573# C a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 VDD B2 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A1 a_940_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X7 a_56_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A2 a_660_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_660_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_2 A1 A2 B1 B2 C VDD VSS ZN
X0 a_1587_96# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X1 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 VSS A2 a_1587_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X3 ZN A1 a_1979_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X4 a_896_96# B1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X5 VSS B2 a_896_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X6 a_504_96# B2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X7 ZN B1 a_504_96# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X8 a_56_573# C a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_244_573# C a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VDD B1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_244_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VDD B2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_1979_96# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X15 ZN A1 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_244_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_56_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_56_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 ZN A2 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi221_4 A1 A2 B1 B2 C VDD VSS ZN
X0 VDD B2 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_1478_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X2 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 a_3320_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X4 ZN A1 a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A1 a_3320_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X6 a_234_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN C VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 a_1822_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN B1 a_662_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X10 VDD B1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_1822_573# C a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_662_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X13 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 a_4136_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X15 a_1822_573# C a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 ZN A2 a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_234_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VSS B2 a_1070_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X19 VSS A2 a_3728_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X20 a_234_573# C a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_1822_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_234_573# C a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_1070_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X24 ZN A2 a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 VDD B2 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 ZN A1 a_1822_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 a_1822_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_1822_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_234_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 a_2912_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X31 VSS A2 a_2912_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X32 VDD B1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 a_3728_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X34 ZN A1 a_4136_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X35 a_244_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X36 VSS C ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X37 ZN B1 a_1478_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
X38 a_234_573# B1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 VSS B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.185u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi221_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 ZN C1 a_291_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS B2 a_827_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_255_573# B1 a_619_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_619_573# B2 a_255_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_255_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD C1 a_255_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A2 a_619_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_619_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_291_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_827_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_1235_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN A1 a_1235_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 VSS C2 a_251_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_2030_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_251_69# C1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_231_573# B1 a_1003_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_1003_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN C1 a_659_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS A2 a_2030_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_231_573# C1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_1003_573# B2 a_231_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN A2 a_1003_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_1191_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN A1 a_1003_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1619_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_231_573# B2 a_1003_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_1003_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD C2 a_231_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 ZN A1 a_2438_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_231_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VDD C1 a_231_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS B2 a_1191_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_659_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 a_1003_573# B1 a_231_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN B1 a_1619_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_2438_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__aoi222_4 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 a_1812_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_652_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN C1 a_652_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_2836_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_1812_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A2 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A1 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS C2 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS B2 a_2010_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_224_573# C1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_4876_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1812_573# A2 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1060_69# C1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 ZN A1 a_4060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD C2 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN A2 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_224_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 ZN C1 a_1468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_1812_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 ZN B1 a_2428_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VSS A2 a_4468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD C1 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_1812_573# B2 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_3244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 ZN B1 a_3244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_224_573# C1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VSS B2 a_2836_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_224_573# B2 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_224_573# B1 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 ZN A1 a_4876_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_1812_573# B1 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VDD C2 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 a_2010_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VSS A2 a_3652_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 a_224_573# B2 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VSS C2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X36 a_3652_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 a_244_69# C1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 a_224_573# B1 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 a_1468_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 a_2428_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 a_224_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X42 a_1812_573# B1 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X43 VDD C1 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X44 a_1812_573# B2 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X45 a_4468_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X46 ZN A1 a_1812_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X47 a_4060_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__aoi222_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_1 I VDD VSS Z
X0 VSS I a_36_146# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 Z a_36_146# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 Z a_36_146# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD I a_36_146# w_n86_453# pmos_6p0 w=0.915u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_2 I VDD VSS Z
X0 VDD I a_36_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VDD a_36_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 Z a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS a_36_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_36_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS I a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_3 I VDD VSS Z
X0 VDD I a_36_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 Z a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD a_36_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_36_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS a_36_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS I a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_36_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_4 I VDD VSS Z
X0 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_8 I VDD VSS Z
X0 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_12 I VDD VSS Z
X0 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_234_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD I a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VSS I a_234_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD I a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_234_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VSS I a_234_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VSS I a_234_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 Z a_234_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_234_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_234_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 a_234_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 VDD a_234_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 VSS a_234_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VDD I a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 Z a_234_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 a_234_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_16 I VDD VSS Z
X0 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X40 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X42 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X44 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X46 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X47 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_20.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__buf_20 I VDD VSS Z
X0 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X36 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X37 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X40 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X42 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X44 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X45 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X46 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X47 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X48 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X49 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X50 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X51 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X52 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X53 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X54 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X55 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X56 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X57 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X58 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X59 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__buf_20.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_1 EN I VDD VSS Z
X0 Z a_468_215# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_468_215# a_36_215# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 Z a_448_693# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD I a_448_693# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X4 VSS EN a_36_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 VDD EN a_36_215# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X6 a_448_693# EN a_468_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 VSS I a_468_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_448_693# EN VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X9 a_468_215# a_36_215# a_448_693# w_n86_453# pmos_6p0 w=0.99u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_2 EN I VDD VSS Z
X0 VDD EN a_38_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 a_450_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X2 VSS a_470_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS I a_470_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_470_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD I a_450_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 Z a_450_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 VDD a_450_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X8 a_450_573# EN a_470_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS EN a_38_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_470_69# a_38_69# a_450_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 a_470_69# a_38_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_3 EN I VDD VSS Z
X0 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_448_573# I VDD w_n86_453# pmos_6p0 w=1.485u l=0.5u
X2 VDD I a_448_573# w_n86_453# pmos_6p0 w=1.485u l=0.5u
X3 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=0.885u l=0.6u
X4 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 Z a_448_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 a_468_69# a_36_69# a_448_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X8 VDD a_448_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 a_448_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_448_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 Z a_448_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=0.885u l=0.6u
X15 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_4 EN I VDD VSS Z
X0 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_448_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X5 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_468_69# a_36_69# a_448_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 VDD I a_448_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 Z a_448_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 a_448_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_448_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 VDD a_448_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X14 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD a_448_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X16 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 Z a_448_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_8 EN I VDD VSS Z
X0 VDD a_428_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X4 a_428_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X5 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_428_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X8 VDD I a_428_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 a_428_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 VDD a_428_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 VDD I a_428_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 Z a_428_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_428_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 VDD a_428_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X16 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 Z a_428_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X18 Z a_428_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_428_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD a_428_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X23 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_468_69# a_36_69# a_428_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X28 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_12 EN I VDD VSS Z
X0 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X4 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X5 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X17 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_476_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X21 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X23 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X24 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X27 a_476_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X30 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X33 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X35 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X36 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 a_468_69# a_36_69# a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X38 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X39 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X41 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__bufz_16 EN I VDD VSS Z
X0 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X17 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X21 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X22 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X23 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X25 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X27 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X28 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X29 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_476_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X32 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X33 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X35 Z a_476_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X36 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X37 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 a_476_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 VDD I a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X41 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X42 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VDD a_476_573# Z w_n86_453# pmos_6p0 w=1.8u l=0.5u
X44 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X46 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X47 VSS I a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X48 VSS a_468_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X49 a_476_573# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X50 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X51 a_468_69# a_36_69# a_476_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X52 a_468_69# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X53 Z a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__bufz_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_1 I VDD VSS Z
X0 Z a_36_140# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X1 VSS I a_36_140# & Metric 1.00 nmos_6p0 w=0.365u l=0.6u
X2 Z a_36_140# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD I a_36_140# w_n86_453# pmos_6p0 w=0.915u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_2 I VDD VSS Z
X0 Z a_36_173# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_36_173# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X2 VDD I a_36_173# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_36_173# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X4 VSS I a_36_173# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 VDD a_36_173# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_3 I VDD VSS Z
X0 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.375u l=0.5u
X1 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.375u l=0.5u
X2 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.6u l=0.6u
X3 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.375u l=0.5u
X4 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.6u l=0.6u
X5 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.55u l=0.6u
X6 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.6u l=0.6u
X7 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.375u l=0.5u
X8 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.375u l=0.5u
X9 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.375u l=0.5u
X10 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.55u l=0.6u
X11 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.6u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_4 I VDD VSS Z
X0 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X1 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X4 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X5 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X7 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X11 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_8 I VDD VSS Z
X0 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X3 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X7 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X8 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X11 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X12 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X15 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X18 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X20 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X23 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_12 I VDD VSS Z
X0 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_268_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X2 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X3 VDD I a_268_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X6 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_268_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS I a_268_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X10 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X11 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X12 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VDD I a_268_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_268_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X16 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X18 a_268_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS I a_268_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X21 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X22 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_268_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X24 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X25 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X28 VDD a_268_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_268_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 VDD I a_268_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X32 Z a_268_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X33 Z a_268_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 VSS I a_268_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X35 VSS a_268_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_16 I VDD VSS Z
X0 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X2 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X7 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X9 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X12 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X14 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X15 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X16 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X19 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X23 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X26 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X29 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X30 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X32 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X33 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X34 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X35 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X37 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X38 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X40 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X41 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X42 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X43 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X44 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X45 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X46 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X47 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_20.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkbuf_20 I VDD VSS Z
X0 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X2 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X7 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X9 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X13 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X15 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X18 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X19 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X21 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X22 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X25 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X28 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X31 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X36 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X37 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X38 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X40 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X41 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X42 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X43 a_224_573# I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X44 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X45 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X46 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X47 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X48 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X49 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X50 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X51 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X52 a_224_573# I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X53 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X54 VSS I a_224_573# & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X55 VDD I a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X56 Z a_224_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X57 VSS a_224_573# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X58 VDD a_224_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X59 Z a_224_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkbuf_20.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_1 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_2 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X3 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_3 I VDD VSS ZN
X0 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X4 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_4 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X3 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X6 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_8 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X3 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X6 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X8 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X10 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X12 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X15 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_12 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X3 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X4 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X6 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X7 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X8 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X11 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X14 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X16 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X17 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X18 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X22 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_16 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X3 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X4 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X8 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X9 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X10 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X14 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X15 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X18 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X20 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X21 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X22 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X24 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X29 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_20.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__clkinv_20 I VDD VSS ZN
X0 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X1 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X2 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X4 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X5 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X7 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X11 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X12 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X13 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X17 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X18 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X19 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X21 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X23 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X25 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X26 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X28 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X30 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X36 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X37 VSS I ZN & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
X38 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 ZN I VSS & Metric 1.00 nmos_6p0 w=0.73u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__clkinv_20.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_1 CLKN D Q VDD VSS
X0 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_1060_156# a_36_175# a_836_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 a_1284_156# a_36_175# a_1060_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 a_1968_592# a_36_175# a_1332_112# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_1264_592# a_448_573# a_1060_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_1332_112# a_1060_156# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VSS a_2360_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_2212_215# a_36_175# a_1968_592# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_1060_156# a_448_573# a_836_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 VDD a_2360_131# a_2212_215# w_n86_453# pmos_6p0 w=1.1u l=0.5u
X10 a_836_156# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_1332_112# a_1264_592# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_2212_215# a_448_573# a_1968_592# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 VSS a_2360_131# a_2212_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X15 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 a_2360_131# a_1968_592# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X17 a_1332_112# a_1060_156# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X19 a_2360_131# a_1968_592# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_836_156# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 VDD a_2360_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_1968_592# a_448_573# a_1332_112# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VSS a_1332_112# a_1284_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_2 CLKN D Q VDD VSS
X0 VDD CLKN a_74_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X1 a_1368_593# a_506_175# a_1078_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VDD a_2412_25# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_506_175# a_74_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X4 a_2272_215# a_74_175# a_1964_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 VSS a_2412_25# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1436_124# a_1078_593# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 a_506_175# a_74_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 a_1078_593# a_506_175# a_874_168# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_2272_215# a_506_175# a_1964_593# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 VDD a_1436_124# a_1368_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_1436_124# a_1078_593# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X12 Q a_2412_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_874_168# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_1964_593# a_506_175# a_1436_124# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 VDD a_2412_25# a_2272_215# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_1078_593# a_74_175# a_874_168# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_2412_25# a_1964_593# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_2412_25# a_1964_593# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS CLKN a_74_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 VSS a_1436_124# a_1388_168# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 a_874_168# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_1388_168# a_74_175# a_1078_593# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X23 VSS a_2412_25# a_2272_215# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 Q a_2412_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_1964_593# a_74_175# a_1436_124# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnq_4 CLKN D Q VDD VSS
X0 a_1981_573# a_474_573# a_1358_115# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 Q a_2412_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS a_2412_25# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD a_1358_115# a_1290_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_1358_115# a_1086_159# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 VSS a_2412_25# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD CLKN a_62_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 VDD a_2412_25# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_474_573# a_62_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 Q a_2412_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_474_573# a_62_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 a_2226_215# a_474_573# a_1981_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X12 a_862_159# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 Q a_2412_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD a_2412_25# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 Q a_2412_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VSS a_1358_115# a_1310_159# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X17 VDD a_2412_25# a_2226_215# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_1086_159# a_62_175# a_862_159# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 VSS CLKN a_62_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_2412_25# a_1981_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_1310_159# a_62_175# a_1086_159# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_2412_25# a_1981_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_1358_115# a_1086_159# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_1981_573# a_62_175# a_1358_115# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_1290_573# a_474_573# a_1086_159# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_2226_215# a_62_175# a_1981_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_1086_159# a_474_573# a_862_159# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 VSS a_2412_25# a_2226_215# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 a_862_159# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1 CLKN D Q RN VDD VSS
X0 a_2799_175# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_1284_175# a_36_175# a_988_573# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X3 a_784_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_2455_131# a_2123_175# a_2799_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_988_573# a_36_175# a_784_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD a_2455_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1296_513# a_988_573# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 a_1192_573# a_436_573# a_988_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_988_573# a_436_573# a_784_573# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 VSS a_2455_131# a_2351_175# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 VDD a_1296_513# a_1192_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 a_2123_175# a_36_175# a_1296_513# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 VSS a_2455_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD a_2455_131# a_2351_175# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_2455_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 a_436_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X18 a_436_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X19 VSS RN a_1452_175# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VDD a_2123_175# a_2455_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_2123_175# a_436_573# a_1296_513# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 a_2351_175# a_436_573# a_2123_175# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X23 a_1192_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_784_573# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X25 a_2351_175# a_36_175# a_2123_175# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_1452_175# a_1296_513# a_1284_175# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X27 a_1296_513# a_988_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2 CLKN D Q RN VDD VSS
X0 VDD a_1332_148# a_1228_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 Q a_2532_392# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS a_2532_392# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1228_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X4 VDD a_2532_392# a_2413_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 VDD a_2532_392# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_2532_392# a_2413_652# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X7 a_820_573# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 a_1452_192# a_1332_148# a_1284_192# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X9 a_1332_148# a_1024_573# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 VSS RN a_1452_192# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 a_2188_652# a_448_573# a_1332_148# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_2413_652# a_36_150# a_2188_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_1284_192# a_36_150# a_1024_573# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 a_448_573# a_36_150# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 a_2413_652# a_448_573# a_2188_652# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X16 a_1332_148# a_1024_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X17 VDD CLKN a_36_150# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_820_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_2188_652# a_36_150# a_1332_148# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 a_2880_192# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X21 a_448_573# a_36_150# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_1024_573# a_36_150# a_820_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 a_1024_573# a_448_573# a_820_573# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 VDD a_2188_652# a_2532_392# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_2532_392# a_2188_652# a_2880_192# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VSS CLKN a_36_150# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X27 Q a_2532_392# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 a_1228_573# a_448_573# a_1024_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 a_2532_392# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4 CLKN D Q RN VDD VSS
X0 a_1332_136# a_1024_593# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_820_593# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 a_2188_640# a_448_573# a_1332_136# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_2413_640# a_36_175# a_2188_640# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 Q a_2532_380# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD a_2532_380# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1284_180# a_36_175# a_1024_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 VSS a_2532_380# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_1024_593# a_36_175# a_820_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 VDD a_2532_380# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_2413_640# a_448_573# a_2188_640# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X12 a_1332_136# a_1024_593# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X13 Q a_2532_380# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS a_2532_380# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_1228_593# a_448_573# a_1024_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_2188_640# a_36_175# a_1332_136# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 a_2880_180# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 VDD a_1332_136# a_1228_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_1024_593# a_448_573# a_820_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VSS RN a_1452_180# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X21 a_1228_593# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X22 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X24 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X25 VDD a_2532_380# a_2413_640# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 VSS a_2532_380# a_2413_640# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X27 VDD a_2188_640# a_2532_380# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_820_593# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X29 Q a_2532_380# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_1452_180# a_1332_136# a_1284_180# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X31 a_2532_380# a_2188_640# a_2880_180# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 Q a_2532_380# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 a_2532_380# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1 CLKN D Q RN SETN VDD VSS
X0 a_1528_215# a_1348_513# a_1360_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_2480_215# a_36_175# a_1348_513# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 a_1360_215# a_36_175# a_1040_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 VSS a_3240_131# a_3192_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_3192_175# SETN a_2704_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 VDD a_1040_573# a_1348_513# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_836_215# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 VSS a_3240_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_1348_513# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X10 VDD a_3240_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_836_215# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_1040_573# a_36_175# a_836_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_1348_513# SETN a_2088_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 a_3240_131# a_2480_215# a_3584_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 a_2480_215# a_448_573# a_1348_513# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_1040_573# a_448_573# a_836_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X17 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 a_2704_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 a_2704_215# a_36_175# a_2480_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X21 a_2704_215# a_448_573# a_2480_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_1244_573# a_448_573# a_1040_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VDD a_3240_131# a_2704_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X24 a_3584_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X25 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 VDD a_1348_513# a_1244_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_3240_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X28 a_1244_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X29 VDD a_2480_215# a_3240_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X30 VSS RN a_1528_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X31 a_2088_215# a_1040_573# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2 CLKN D Q RN SETN VDD VSS
X0 VDD a_1379_171# a_1225_589# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VDD a_2437_215# a_3225_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X2 a_1379_171# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_1331_215# a_57_150# a_1021_589# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_3569_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_1225_589# a_469_573# a_1021_589# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_2437_215# a_469_573# a_1379_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_1021_589# a_469_573# a_817_589# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_2661_215# a_469_573# a_2437_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_469_573# a_57_150# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_2661_215# a_57_150# a_2437_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD CLKN a_57_150# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_469_573# a_57_150# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 VSS RN a_1499_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 a_2045_215# a_1021_589# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 VSS a_3225_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 Q a_3225_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 Q a_3225_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VSS a_3225_131# a_3161_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 a_817_589# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X20 a_1225_589# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X21 VSS CLKN a_57_150# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_2437_215# a_57_150# a_1379_171# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X23 VDD a_3225_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VDD a_1021_589# a_1379_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_2661_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 a_1499_215# a_1379_171# a_1331_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_1379_171# SETN a_2045_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 VDD a_3225_131# a_2661_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X29 a_817_589# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_3225_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X31 a_3161_175# SETN a_2661_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X32 a_1021_589# a_57_150# a_817_589# w_n86_453# pmos_6p0 w=1u l=0.5u
X33 a_3225_131# a_2437_215# a_3569_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4 CLKN D Q RN SETN VDD VSS
X0 VDD a_3209_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 Q a_3209_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_1020_573# a_36_175# a_816_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 VDD a_1332_171# a_1224_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 VDD a_3209_131# a_2676_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 a_2060_215# a_1020_573# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 a_3209_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 a_3209_131# a_2452_215# a_3553_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 VDD a_1020_573# a_1332_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 Q a_3209_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD a_2452_215# a_3209_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_2452_215# a_36_175# a_1332_171# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 a_1224_573# a_448_573# a_1020_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_3553_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 a_816_573# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 VSS a_3209_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_1452_215# a_1332_171# a_1284_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 VSS a_3209_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VDD a_3209_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 a_1332_171# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X21 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 a_1284_215# a_36_175# a_1020_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_1332_171# SETN a_2060_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 Q a_3209_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_2452_215# a_448_573# a_1332_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_1224_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 Q a_3209_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X30 VSS a_3209_131# a_3161_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X31 a_2676_215# a_36_175# a_2452_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_2676_215# a_448_573# a_2452_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X33 VSS RN a_1452_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X34 a_2676_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X35 a_3161_175# SETN a_2676_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X36 a_1020_573# a_448_573# a_816_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X37 a_816_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnrsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1 CLKN D Q SETN VDD VSS
X0 VDD a_1276_425# a_1228_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_820_573# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 VDD CLKN a_36_146# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 VSS a_1276_425# a_1288_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_1688_215# a_1024_573# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 a_3076_171# a_2080_215# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X6 a_428_573# a_36_146# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 a_2340_183# a_36_146# a_2080_215# w_n86_453# pmos_6p0 w=1.1u l=0.5u
X8 VSS CLKN a_36_146# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 a_1288_215# a_36_146# a_1024_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 VDD SETN a_1276_425# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_2936_183# SETN a_2340_183# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X12 VDD a_3076_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_2080_215# a_36_146# a_1276_425# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 VSS a_3076_171# a_2936_183# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 a_820_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VSS a_3076_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_1024_573# a_428_573# a_820_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 VDD a_3076_171# a_2340_183# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_3076_171# a_2080_215# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X20 a_1024_573# a_36_146# a_820_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X21 a_1276_425# a_1024_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X22 a_2340_183# a_428_573# a_2080_215# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X23 a_2080_215# a_428_573# a_1276_425# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_428_573# a_36_146# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X25 a_2340_183# SETN VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X26 a_1228_573# a_428_573# a_1024_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_1276_425# SETN a_1688_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2 CLKN D Q SETN VDD VSS
X0 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_3064_171# a_2068_195# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X2 VSS a_3064_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_836_195# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_2328_163# a_36_175# a_2068_195# w_n86_453# pmos_6p0 w=1.1u l=0.5u
X5 VDD a_3064_171# a_2328_163# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_1040_586# a_36_175# a_836_195# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_836_195# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 VSS a_1332_151# a_1284_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_2068_195# a_36_175# a_1332_151# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 a_2924_183# SETN a_2328_163# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X11 a_3064_171# a_2068_195# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X12 a_2068_195# a_448_573# a_1332_151# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_2328_163# a_448_573# a_2068_195# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X14 VSS a_3064_171# a_2924_183# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 Q a_3064_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1284_195# a_36_175# a_1040_586# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X17 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 VDD SETN a_1332_151# w_n86_453# pmos_6p0 w=1u l=0.5u
X20 Q a_3064_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_1332_151# SETN a_1676_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 VDD a_1332_151# a_1264_586# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 VDD a_3064_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_1040_586# a_448_573# a_836_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X26 a_1332_151# a_1040_586# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_2328_163# SETN VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X28 a_1676_195# a_1040_586# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_1264_586# a_448_573# a_1040_586# w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4 CLKN D Q SETN VDD VSS
X0 VSS CLKN a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 VDD a_3156_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_840_215# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 Q a_3156_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_2420_183# a_448_573# a_2160_215# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X5 a_2420_183# SETN VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X6 Q a_3156_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1044_582# a_448_573# a_840_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_2160_215# a_448_573# a_1296_425# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_1296_425# SETN a_1708_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 Q a_3156_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_1296_425# a_1044_582# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X12 VDD a_3156_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 Q a_3156_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 a_3016_183# SETN a_2420_183# & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X15 a_3156_171# a_2160_215# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X16 a_840_215# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_2420_183# a_36_175# a_2160_215# w_n86_453# pmos_6p0 w=1.1u l=0.5u
X18 a_2160_215# a_36_175# a_1296_425# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 VDD a_3156_171# a_2420_183# w_n86_453# pmos_6p0 w=1u l=0.5u
X20 a_3156_171# a_2160_215# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X21 a_1044_582# a_36_175# a_840_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 VDD CLKN a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X24 VSS a_1296_425# a_1308_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_1708_215# a_1044_582# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X26 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X27 VSS a_3156_171# a_3016_183# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_1248_582# a_448_573# a_1044_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 a_1308_215# a_36_175# a_1044_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X30 VDD a_1296_425# a_1248_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X31 VDD SETN a_1296_425# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 VSS a_3156_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VSS a_3156_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffnsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_1 CLK D Q VDD VSS
X0 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_1820_573# a_448_573# a_1276_173# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 a_836_217# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X3 VSS a_1276_173# a_1228_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X4 a_1264_573# a_36_175# a_1004_217# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_1276_173# a_1004_217# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X6 a_2192_173# a_1820_573# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X7 a_1004_217# D a_856_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_2144_217# a_36_175# a_1820_573# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X9 VDD a_1276_173# a_1264_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_2160_573# a_448_573# a_1820_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_1228_217# a_448_573# a_1004_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X12 VDD a_2192_173# a_2160_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 Q a_2192_173# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 a_1004_217# D a_836_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X17 a_1276_173# a_1004_217# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_1820_573# a_36_175# a_1276_173# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 a_2192_173# a_1820_573# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X21 Q a_2192_173# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_856_573# a_448_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VSS a_2192_173# a_2144_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_2 CLK D Q VDD VSS
X0 VSS a_1318_171# a_1270_215# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X1 a_1942_582# a_448_573# a_1318_171# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 VSS a_2234_172# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 Q a_2234_172# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD CLK a_36_146# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_2234_172# a_1942_582# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1270_215# a_448_573# a_1046_215# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X7 VSS a_2234_172# a_2186_216# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X8 VDD a_2234_172# a_2202_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 VSS CLK a_36_146# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_1318_171# a_1046_215# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_2186_216# a_36_146# a_1942_582# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X12 a_2234_172# a_1942_582# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_1318_171# a_1046_215# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X14 a_2202_582# a_448_573# a_1942_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 a_1046_215# D a_878_215# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X16 a_1270_582# a_36_146# a_1046_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_898_582# a_448_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_1942_582# a_36_146# a_1318_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_878_215# a_36_146# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X20 a_448_573# a_36_146# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 VDD a_2234_172# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 Q a_2234_172# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_448_573# a_36_146# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X24 a_1046_215# D a_898_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 VDD a_1318_171# a_1270_582# w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffq_4 CLK D Q VDD VSS
X0 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_1899_573# a_448_573# a_1276_173# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 a_836_217# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X3 a_1276_173# a_1004_217# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X4 VSS a_1276_173# a_1228_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X5 a_1276_173# a_1004_217# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X6 a_1004_217# D a_856_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_2192_173# a_1899_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 Q a_2192_173# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD a_1899_573# a_2192_173# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_2144_217# a_36_175# a_1899_573# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X11 a_1248_573# a_36_175# a_1004_217# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 VDD a_2192_173# a_2184_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 Q a_2192_173# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 Q a_2192_173# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD a_1276_173# a_1248_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_1899_573# a_36_175# a_1276_173# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 VDD a_2192_173# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_1228_217# a_448_573# a_1004_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X19 VSS a_1899_573# a_2192_173# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_1004_217# D a_836_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X23 Q a_2192_173# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VSS a_2192_173# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 a_2184_573# a_448_573# a_1899_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 VSS a_2192_173# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 VDD a_2192_173# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_2192_173# a_1899_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_856_573# a_448_573# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X31 VSS a_2192_173# a_2144_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_1 CLK D Q RN VDD VSS
X0 a_1232_593# a_40_175# a_1028_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_2160_170# a_40_175# a_1336_126# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VDD a_2160_170# a_2488_126# w_n86_453# pmos_6p0 w=0.98u l=0.5u
X3 VSS RN a_1456_170# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 VDD a_1336_126# a_1232_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_1288_170# a_432_573# a_1028_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 a_2384_170# a_432_573# a_2160_170# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_2488_126# a_2160_170# a_2832_170# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 a_1232_593# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_1336_126# a_1028_593# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_2160_170# a_432_573# a_1336_126# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 a_2832_170# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X12 a_432_573# a_40_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X13 a_1028_593# a_40_175# a_824_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 VSS a_2488_126# a_2384_170# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 VDD a_2488_126# a_2384_170# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VSS a_2488_126# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD a_2488_126# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_824_593# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X19 VSS CLK a_40_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_824_593# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X21 a_1028_593# a_432_573# a_824_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 VDD CLK a_40_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_2384_170# a_40_175# a_2160_170# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 a_432_573# a_40_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X25 a_1456_170# a_1336_126# a_1288_170# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X26 a_1336_126# a_1028_593# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X27 a_2488_126# RN VDD w_n86_453# pmos_6p0 w=0.98u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_2 CLK D Q RN VDD VSS
X0 a_820_593# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_1024_593# a_36_170# a_820_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 VSS a_2478_125# a_2374_169# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X3 a_1024_593# a_448_573# a_820_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_1332_125# a_1024_593# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X5 a_2478_125# a_2150_169# a_2822_169# & Metric 1.00 nmos_6p0 w=1.18u l=0.6u
X6 a_1228_593# a_36_170# a_1024_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VSS CLK a_36_170# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 VDD a_1332_125# a_1228_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_2150_169# a_36_170# a_1332_125# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 Q a_2478_125# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_2374_169# a_448_573# a_2150_169# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_2374_169# a_36_170# a_2150_169# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_1228_593# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_1332_125# a_1024_593# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X15 VDD a_2478_125# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_820_593# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 VSS a_2478_125# Q & Metric 1.00 nmos_6p0 w=1.25u l=0.6u
X18 VDD a_2478_125# a_2374_169# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_1452_169# a_1332_125# a_1284_169# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VDD CLK a_36_170# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_2478_125# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 VSS RN a_1452_169# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X23 a_448_573# a_36_170# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X24 a_1284_169# a_448_573# a_1024_593# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X25 VDD a_2150_169# a_2478_125# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 Q a_2478_125# VSS & Metric 1.00 nmos_6p0 w=1.25u l=0.6u
X27 a_2150_169# a_448_573# a_1332_125# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X28 a_2822_169# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X29 a_448_573# a_36_170# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrnq_4 CLK D Q RN VDD VSS
X0 Q a_2473_160# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_796_582# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 VSS a_2473_160# a_2369_204# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_1204_582# a_36_175# a_1000_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 VDD a_2473_160# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_1456_204# a_1308_538# a_1288_204# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 a_2473_160# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_2473_160# a_2145_204# a_2817_204# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD a_1308_538# a_1204_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_2145_204# a_36_175# a_1308_538# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_2145_204# a_2473_160# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1204_582# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_1288_204# a_448_573# a_1000_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 VSS RN a_1456_204# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 a_2369_204# a_448_573# a_2145_204# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VDD a_2473_160# a_2369_204# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_2369_204# a_36_175# a_2145_204# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 a_796_582# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X19 VSS a_2473_160# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_1000_582# a_36_175# a_796_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X23 a_2817_204# RN VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 VSS a_2473_160# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_1308_538# a_1000_582# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X27 Q a_2473_160# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_2145_204# a_448_573# a_1308_538# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_1000_582# a_448_573# a_796_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_1308_538# a_1000_582# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X31 Q a_2473_160# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 VDD a_2473_160# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 Q a_2473_160# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1 CLK D Q RN SETN VDD VSS
X0 a_2528_215# a_428_586# a_2304_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_3467_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_776_582# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_980_582# a_428_586# a_776_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_776_582# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 VSS RN a_1468_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 VDD a_3123_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1468_215# a_1288_538# a_1300_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 VSS a_3123_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_428_586# a_36_586# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_1184_582# a_36_586# a_980_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_3123_131# a_2528_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_1300_215# a_428_586# a_980_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 VDD a_1288_538# a_1184_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_3123_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X15 VSS a_3123_131# a_3075_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 a_2528_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 VDD a_980_582# a_1288_538# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_1288_538# SETN a_1912_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 a_1288_538# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X20 VDD a_2304_215# a_3123_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_1912_215# a_980_582# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 VSS CLK a_36_586# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 a_980_582# a_36_586# a_776_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_2528_215# a_36_586# a_2304_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_1184_582# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X26 VDD CLK a_36_586# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X27 a_2304_215# a_428_586# a_1288_538# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_3123_131# a_2304_215# a_3467_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X29 a_2304_215# a_36_586# a_1288_538# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_3075_175# SETN a_2528_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X31 a_428_586# a_36_586# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2 CLK D Q RN SETN VDD VSS
X0 a_1184_573# a_36_175# a_980_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_2316_215# a_36_175# a_1288_529# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 VSS a_3132_131# a_3084_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 a_1924_215# a_980_573# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 VDD a_1288_529# a_1184_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_2540_215# a_428_573# a_2316_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 a_776_573# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 VDD a_3132_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS RN a_1468_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X11 VSS a_3132_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_428_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 a_1468_215# a_1288_529# a_1300_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 Q a_3132_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 Q a_3132_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_1300_215# a_428_573# a_980_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X17 VDD a_3132_131# a_2540_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_3132_131# a_2316_215# a_3476_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 a_3084_175# SETN a_2540_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_3132_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_2540_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 VDD a_980_573# a_1288_529# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VDD a_2316_215# a_3132_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X24 a_428_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X25 a_1288_529# SETN a_1924_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X26 a_3476_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X27 a_776_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_980_573# a_36_175# a_776_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_980_573# a_428_573# a_776_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_2540_215# a_36_175# a_2316_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X31 a_1184_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_1288_529# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X33 a_2316_215# a_428_573# a_1288_529# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4 CLK D Q RN SETN VDD VSS
X0 a_1184_573# a_36_175# a_980_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_2316_215# a_36_175# a_1288_529# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 VSS a_3132_131# a_3084_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 Q a_3132_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_1924_215# a_980_573# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 VDD a_1288_529# a_1184_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_2540_215# a_428_573# a_2316_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X9 a_776_573# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 Q a_3132_131# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD a_3132_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS RN a_1468_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 a_428_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_1468_215# a_1288_529# a_1300_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 Q a_3132_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 Q a_3132_131# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VDD a_3132_131# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_1300_215# a_428_573# a_980_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 VDD a_3132_131# a_2540_215# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 a_3132_131# a_2316_215# a_3476_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X21 a_3084_175# SETN a_2540_215# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_3132_131# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_2540_215# SETN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X24 VDD a_980_573# a_1288_529# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 VDD a_2316_215# a_3132_131# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 a_428_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X27 a_1288_529# SETN a_1924_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_3476_175# RN VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X29 a_776_573# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_980_573# a_36_175# a_776_573# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X31 a_980_573# a_428_573# a_776_573# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_2540_215# a_36_175# a_2316_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X33 a_1184_573# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X34 VSS a_3132_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X35 a_1288_529# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X36 a_2316_215# a_428_573# a_1288_529# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X37 VSS a_3132_131# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffrsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_1 CLK D Q SETN VDD VSS
X0 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 VSS a_3056_171# a_2992_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 a_3056_171# a_2152_215# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X3 a_2152_215# a_448_573# a_1332_135# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_1332_135# a_1060_179# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_1744_215# a_1060_179# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 a_836_179# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 VDD SETN a_1332_135# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_2152_215# a_36_175# a_1332_135# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 VSS a_1332_135# a_1284_179# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 a_1060_179# a_448_573# a_836_179# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_1332_135# a_1264_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_1284_179# a_448_573# a_1060_179# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 VDD a_3056_171# a_2376_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 Q a_3056_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_1264_593# a_36_175# a_1060_179# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X18 a_2376_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_2992_215# SETN a_2376_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X20 a_2376_215# a_36_175# a_2152_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_1060_179# a_36_175# a_836_179# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X23 a_1332_135# SETN a_1744_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_3056_171# a_2152_215# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X25 a_2376_215# a_448_573# a_2152_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_836_179# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 Q a_3056_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_2 CLK D Q SETN VDD VSS
X0 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_2350_215# a_448_573# a_2126_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 Q a_3030_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD a_3030_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_2350_215# a_36_175# a_2126_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 a_1346_150# a_1060_194# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_1296_194# a_448_573# a_1060_194# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 VSS a_3030_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD a_1346_150# a_1293_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_3030_171# a_2126_215# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_3030_171# a_2126_215# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS a_1346_150# a_1296_194# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X12 a_1734_215# a_1060_194# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 a_1060_194# a_36_175# a_836_194# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 a_1060_194# a_448_573# a_836_194# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 VSS a_3030_171# a_2982_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 VDD a_3030_171# a_2350_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_2126_215# a_448_573# a_1346_150# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X19 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_1293_593# a_36_175# a_1060_194# w_n86_453# pmos_6p0 w=1u l=0.5u
X21 VDD SETN a_1346_150# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 a_2126_215# a_36_175# a_1346_150# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X24 a_2350_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X25 Q a_3030_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_836_194# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_836_194# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_2982_215# SETN a_2350_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_1346_150# SETN a_1734_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dffsnq_4 CLK D Q SETN VDD VSS
X0 VSS CLK a_36_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 VSS a_3017_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_3017_171# a_2113_215# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS a_1353_171# a_1284_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 Q a_3017_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD a_2113_215# a_3017_171# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_3017_171# a_2969_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 Q a_3017_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_3017_171# a_2113_215# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_1353_171# SETN a_1697_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 a_2113_215# a_448_573# a_1353_171# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X11 VDD a_3017_171# a_2337_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_836_215# D VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 VDD a_3017_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 Q a_3017_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_2337_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_1060_215# a_448_573# a_836_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_2113_215# a_36_175# a_1353_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 Q a_3017_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VDD a_1353_171# a_1293_593# w_n86_453# pmos_6p0 w=1u l=0.5u
X20 VDD a_3017_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VDD CLK a_36_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_448_573# a_36_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 a_1284_215# a_448_573# a_1060_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_1293_593# a_36_175# a_1060_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_1353_171# a_1060_215# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_1697_215# a_1060_215# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_2969_215# SETN a_2337_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_448_573# a_36_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X29 VDD SETN a_1353_171# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_2337_215# a_448_573# a_2113_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X31 a_836_215# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_2337_215# a_36_175# a_2113_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X33 VSS a_3017_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 a_1060_215# a_36_175# a_836_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X35 VSS a_2113_215# a_3017_171# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dffsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_1 I VDD VSS Z
X0 VSS I a_36_254# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X1 Z a_598_123# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS a_448_646# a_598_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 a_448_646# a_36_254# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X4 Z a_598_123# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_448_646# a_36_254# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 VDD I a_36_254# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X7 VDD a_448_646# a_598_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_2 I VDD VSS Z
X0 VSS a_589_123# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VDD a_448_695# a_589_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X2 Z a_589_123# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_448_695# a_36_259# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X4 a_448_695# a_36_259# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_448_695# a_589_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 VSS I a_36_259# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X7 VDD I a_36_259# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X8 VDD a_589_123# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 Z a_589_123# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlya_4 I VDD VSS Z
X0 Z a_629_152# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_629_152# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD a_629_152# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD a_449_686# a_629_152# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X4 Z a_629_152# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 Z a_629_152# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_449_686# a_37_152# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X7 a_449_686# a_37_152# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 Z a_629_152# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS a_629_152# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VSS a_449_686# a_629_152# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 VDD a_629_152# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VDD I a_37_152# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X13 VSS I a_37_152# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlya_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_1 I VDD VSS Z
X0 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 a_506_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X2 a_486_658# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X3 VDD a_298_267# a_698_662# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X4 a_486_658# a_36_123# a_298_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_298_267# a_698_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 a_918_662# a_298_267# a_698_662# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X7 Z a_918_662# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_918_662# a_298_267# a_698_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X10 Z a_918_662# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_506_123# a_36_123# a_298_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_2 I VDD VSS Z
X0 Z a_918_637# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_918_637# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_506_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 a_918_637# a_298_267# a_698_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X4 VDD a_298_267# a_698_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X6 VDD a_918_637# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_486_637# a_36_123# a_298_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X8 VSS a_298_267# a_698_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 a_918_637# a_298_267# a_698_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X10 a_486_637# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X11 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 Z a_918_637# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_506_123# a_36_123# a_298_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyb_4 I VDD VSS Z
X0 Z a_929_666# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_517_123# a_47_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X2 VSS a_929_666# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_497_666# a_47_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X4 VSS a_929_666# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_497_666# a_47_123# a_309_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X6 VDD a_929_666# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 Z a_929_666# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_929_666# a_309_267# a_709_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 VSS I a_47_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X10 VSS a_309_267# a_709_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 VDD a_309_267# a_709_666# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X12 a_517_123# a_47_123# a_309_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X13 Z a_929_666# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_929_666# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD a_929_666# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD I a_47_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X17 a_929_666# a_309_267# a_709_666# w_n86_453# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyb_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_1 I VDD VSS Z
X0 a_497_630# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 a_517_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X2 a_497_630# a_36_123# a_309_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X3 Z a_1729_630# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_929_630# a_309_267# a_709_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X5 VDD a_1109_212# a_1509_630# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X6 a_1317_68# a_929_630# a_1109_212# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X7 a_1729_630# a_1109_212# a_1509_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 VSS a_309_267# a_709_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 a_1729_630# a_1109_212# a_1509_630# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X10 VDD a_309_267# a_709_630# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X11 VSS a_1109_212# a_1509_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 a_1297_630# a_929_630# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X13 a_929_630# a_309_267# a_709_630# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X14 a_517_123# a_36_123# a_309_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X15 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X16 a_1297_630# a_929_630# a_1109_212# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X17 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X18 a_1317_68# a_929_630# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X19 Z a_1729_630# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_2 I VDD VSS Z
X0 a_1718_637# a_1098_212# a_1498_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 VDD a_1098_212# a_1498_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X2 a_506_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 VSS a_1718_637# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_918_637# a_298_267# a_698_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_298_267# a_698_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 a_1286_637# a_918_637# a_1098_212# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X7 VDD a_298_267# a_698_637# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X8 a_918_637# a_298_267# a_698_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 a_1286_637# a_918_637# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X10 a_1306_68# a_918_637# a_1098_212# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 a_1718_637# a_1098_212# a_1498_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 VSS a_1098_212# a_1498_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X13 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X14 Z a_1718_637# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_486_637# a_36_123# a_298_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X16 a_486_637# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X17 a_1306_68# a_918_637# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X18 Z a_1718_637# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X20 a_506_123# a_36_123# a_298_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X21 VDD a_1718_637# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyc_4 I VDD VSS Z
X0 a_1272_596# a_904_596# a_1084_261# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 Z a_1704_596# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_1292_117# a_904_596# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 a_904_596# a_284_284# a_684_117# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X4 a_1292_117# a_904_596# a_1084_261# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X5 a_472_596# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X6 VDD a_1704_596# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_472_596# a_36_123# a_284_284# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X8 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X9 VDD a_1084_261# a_1484_596# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X10 VDD a_1704_596# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS a_1704_596# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_1704_596# a_1084_261# a_1484_596# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X13 a_492_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X14 VSS a_1084_261# a_1484_117# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X15 VSS a_1704_596# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1704_596# a_1084_261# a_1484_117# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X17 Z a_1704_596# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 Z a_1704_596# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VDD a_284_284# a_684_596# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X20 a_492_123# a_36_123# a_284_284# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X21 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X22 a_1272_596# a_904_596# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X23 Z a_1704_596# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_904_596# a_284_284# a_684_596# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X25 VSS a_284_284# a_684_117# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyc_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_1 I VDD VSS Z
X0 a_2107_116# a_1719_633# a_1899_260# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X1 VDD I a_37_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X2 VSS I a_37_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 a_1719_633# a_1099_260# a_1499_116# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X4 a_919_633# a_299_267# a_699_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VDD a_1899_260# a_2300_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X6 a_507_123# a_37_123# a_299_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X7 a_1287_633# a_919_633# a_1099_260# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X8 Z a_2520_633# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_487_633# a_37_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X10 a_507_123# a_37_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 VSS a_299_267# a_699_116# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 a_2520_633# a_1899_260# a_2300_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X13 a_1307_116# a_919_633# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X14 a_919_633# a_299_267# a_699_116# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X15 a_1307_116# a_919_633# a_1099_260# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X16 a_487_633# a_37_123# a_299_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X17 a_2087_633# a_1719_633# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X18 VDD a_1099_260# a_1499_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X19 a_2087_633# a_1719_633# a_1899_260# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X20 a_2520_633# a_1899_260# a_2300_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X21 a_1719_633# a_1099_260# a_1499_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X22 VSS a_1899_260# a_2300_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X23 a_2107_116# a_1719_633# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X24 VDD a_299_267# a_699_633# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X25 a_1287_633# a_919_633# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X26 Z a_2520_633# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VSS a_1099_260# a_1499_116# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_2 I VDD VSS Z
X0 a_1286_639# a_918_639# a_1098_212# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 a_2518_639# a_1898_258# a_2298_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X2 Z a_2518_639# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_2106_114# a_1718_639# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X4 VDD a_298_267# a_698_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_1098_212# a_1498_114# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 a_1286_639# a_918_639# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X7 a_506_123# a_36_123# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 VDD a_1898_258# a_2298_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X9 VDD I a_36_123# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X10 VSS a_298_267# a_698_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 a_486_639# a_36_123# a_298_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X12 a_486_639# a_36_123# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X13 a_918_639# a_298_267# a_698_68# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X14 a_1306_68# a_918_639# a_1098_212# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X15 VSS a_2518_639# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD a_2518_639# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_2086_639# a_1718_639# a_1898_258# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X18 a_1718_639# a_1098_212# a_1498_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X19 VSS a_1898_258# a_2298_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X20 a_2086_639# a_1718_639# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X21 VDD a_1098_212# a_1498_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X22 a_1306_68# a_918_639# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X23 a_2518_639# a_1898_258# a_2298_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X24 VSS I a_36_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X25 a_2106_114# a_1718_639# a_1898_258# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X26 a_506_123# a_36_123# a_298_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X27 a_1718_639# a_1098_212# a_1498_114# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X28 a_918_639# a_298_267# a_698_639# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X29 Z a_2518_639# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__dlyd_4 I VDD VSS Z
X0 a_1288_640# a_920_640# a_1100_268# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X1 VDD a_2520_640# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_2520_640# a_1900_267# a_2300_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X3 Z a_2520_640# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_488_640# a_38_124# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X5 VSS a_1900_267# a_2300_69# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 a_920_640# a_300_268# a_700_124# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X7 Z a_2520_640# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_488_640# a_38_124# a_300_268# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X9 a_1308_124# a_920_640# a_1100_268# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X10 VSS a_2520_640# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS a_300_268# a_700_124# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 VSS a_2520_640# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD a_1100_268# a_1500_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X14 a_2088_640# a_1720_640# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X15 a_1308_124# a_920_640# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X16 Z a_2520_640# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VSS I a_38_124# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X18 a_1720_640# a_1100_268# a_1500_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X19 a_2108_123# a_1720_640# a_1900_267# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X20 a_1720_640# a_1100_268# a_1500_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X21 a_2088_640# a_1720_640# a_1900_267# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X22 a_508_124# a_38_124# a_300_268# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X23 VDD a_2520_640# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VDD a_300_268# a_700_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X25 Z a_2520_640# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VSS a_1100_268# a_1500_123# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X27 a_2108_123# a_1720_640# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X28 VDD a_1900_267# a_2300_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X29 a_508_124# a_38_124# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X30 a_1288_640# a_920_640# VDD w_n86_453# pmos_6p0 w=0.36u l=0.5u
X31 VDD I a_38_124# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X32 a_920_640# a_300_268# a_700_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X33 a_2520_640# a_1900_267# a_2300_640# w_n86_453# pmos_6p0 w=0.36u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__dlyd_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__endcap.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__endcap VSS VDD
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__endcap.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_1 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_2 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_4 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_8 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_16 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_32.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_32 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_32.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_64.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fill_64 VDD VSS
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fill_64.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_4 VDD VSS
X0 VDD a_124_481# a_36_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X1 a_124_481# a_36_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_8 VDD VSS
X0 VDD a_124_481# a_36_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X1 VDD a_572_481# a_484_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X2 a_572_481# a_484_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X3 a_124_481# a_36_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_16 VDD VSS
X0 VDD a_1468_481# a_1380_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X1 VDD a_124_481# a_36_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X2 VDD a_572_481# a_484_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X3 a_1020_481# a_932_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X4 a_572_481# a_484_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X5 a_124_481# a_36_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X6 VDD a_1020_481# a_932_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X7 a_1468_481# a_1380_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_32.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_32 VDD VSS
X0 a_2364_481# a_2276_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X1 VDD a_1468_481# a_1380_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X2 a_3260_481# a_3172_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X3 VDD a_124_481# a_36_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X4 VDD a_572_481# a_484_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X5 VDD a_2364_481# a_2276_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X6 VDD a_1916_481# a_1828_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X7 a_1020_481# a_932_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X8 VDD a_3260_481# a_3172_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X9 a_572_481# a_484_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X10 a_124_481# a_36_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X11 VDD a_1020_481# a_932_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X12 VDD a_2812_481# a_2724_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X13 a_1916_481# a_1828_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X14 a_1468_481# a_1380_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X15 a_2812_481# a_2724_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_32.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_64.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__fillcap_64 VDD VSS
X0 VDD a_6396_481# a_6308_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X1 a_2364_481# a_2276_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X2 VDD a_1468_481# a_1380_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X3 VDD a_4156_481# a_4068_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X4 VDD a_5948_481# a_5860_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X5 a_5948_481# a_5860_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X6 a_3260_481# a_3172_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X7 VDD a_124_481# a_36_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X8 VDD a_3708_481# a_3620_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X9 a_6844_481# a_6756_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X10 a_6396_481# a_6308_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X11 VDD a_572_481# a_484_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X12 VDD a_2364_481# a_2276_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X13 VDD a_6844_481# a_6756_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X14 VDD a_5052_481# a_4964_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X15 VDD a_1916_481# a_1828_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X16 a_3708_481# a_3620_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X17 a_1020_481# a_932_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X18 VDD a_4604_481# a_4516_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X19 a_4604_481# a_4516_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X20 a_4156_481# a_4068_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X21 a_5500_481# a_5412_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X22 VDD a_3260_481# a_3172_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X23 a_572_481# a_484_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X24 a_124_481# a_36_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X25 a_5052_481# a_4964_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X26 VDD a_1020_481# a_932_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X27 VDD a_2812_481# a_2724_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X28 a_1916_481# a_1828_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X29 VDD a_5500_481# a_5412_573# w_n86_453# pmos_6p0 w=1.83u l=1u
X30 a_1468_481# a_1380_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
X31 a_2812_481# a_2724_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=1u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__fillcap_64.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__filltie.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__filltie VSS VDD
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__filltie.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__hold.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__hold Z VSS VDD
X0 VDD a_172_123# Z w_n86_453# pmos_6p0 w=0.36u l=2u
X1 VSS a_172_123# Z & Metric 1.00 nmos_6p0 w=0.36u l=2u
X2 a_172_123# Z VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_172_123# Z VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__hold.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_1 CLKN E Q TE VDD VSS
X0 VSS TE a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_1908_573# a_1012_112# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_572_112# a_582_476# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 a_682_576# a_582_476# a_458_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X4 a_682_576# a_572_112# a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X5 a_2628_157# a_1908_573# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 VDD a_682_576# a_1012_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 VSS a_1012_112# a_916_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 Q a_2628_157# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X9 Q a_2628_157# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS CLKN a_582_476# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 a_1908_573# a_1012_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_310_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 VSS a_682_576# a_1012_112# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 a_458_576# E a_310_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X15 a_984_576# a_572_112# a_682_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X16 a_36_156# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 VDD CLKN a_582_476# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_916_156# a_582_476# a_682_576# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X19 VSS CLKN a_2628_157# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 a_2624_573# a_1908_573# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_2628_157# CLKN a_2624_573# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_572_112# a_582_476# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X23 VDD a_1012_112# a_984_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_2 CLKN E Q TE VDD VSS
X0 VSS TE a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_1900_161# a_964_112# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_572_112# a_680_532# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 Q a_2580_161# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_692_156# a_572_112# a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X5 a_462_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X6 VDD a_2580_161# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_2580_161# a_1900_161# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X8 a_2580_161# CLKN a_2580_573# w_n86_453# pmos_6p0 w=1.68u l=0.5u
X9 a_572_112# a_680_532# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 VSS a_2580_161# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X11 a_692_156# a_680_532# a_610_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 VSS a_692_156# a_964_112# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_610_576# E a_462_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_984_576# a_572_112# a_692_156# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X15 VSS a_964_112# a_916_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X16 a_36_156# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 VDD a_692_156# a_964_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 VSS CLKN a_680_532# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X19 a_916_156# a_680_532# a_692_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VDD CLKN a_680_532# w_n86_453# pmos_6p0 w=1.68u l=0.5u
X21 VSS CLKN a_2580_161# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X22 Q a_2580_161# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X23 a_2580_573# a_1900_161# VDD w_n86_453# pmos_6p0 w=1.68u l=0.5u
X24 VDD a_964_112# a_984_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X25 a_1900_161# a_964_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtn_4 CLKN E Q TE VDD VSS
X0 VSS TE a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 Q a_2591_156# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X2 VDD a_695_156# a_967_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 VSS a_2591_156# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X4 a_987_576# a_575_112# a_695_156# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 VDD CLKN a_683_532# w_n86_453# pmos_6p0 w=1.68u l=0.5u
X6 VSS a_967_112# a_919_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X7 a_1891_573# a_967_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 a_2591_156# a_1891_573# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X9 a_2591_585# a_1891_573# VDD w_n86_453# pmos_6p0 w=1.68u l=0.5u
X10 a_919_156# a_683_532# a_695_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 Q a_2591_156# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_440_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 VDD a_2591_156# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS a_695_156# a_967_112# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 a_588_576# E a_440_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X16 Q a_2591_156# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X17 VDD a_967_112# a_987_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_2591_156# CLKN a_2591_585# w_n86_453# pmos_6p0 w=1.68u l=0.5u
X19 Q a_2591_156# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS CLKN a_683_532# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X21 VSS a_2591_156# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X22 a_575_112# a_683_532# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_36_156# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 VDD a_2591_156# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_695_156# a_575_112# a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X26 VSS CLKN a_2591_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X27 a_575_112# a_683_532# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X28 a_695_156# a_683_532# a_588_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X29 a_1891_573# a_967_112# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtn_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_1 CLK E Q TE VDD VSS
X0 a_616_112# CLK VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X1 a_644_576# a_616_112# a_36_137# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_1008_112# a_644_576# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X3 a_616_112# CLK VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 Q a_2207_137# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X5 a_36_137# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 Q a_2207_137# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_344_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 a_492_576# E a_344_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X9 a_644_576# a_544_476# a_492_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X10 a_1028_576# a_616_112# a_644_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 a_2207_137# CLK VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 VSS a_616_112# a_544_476# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 VSS a_1008_112# a_960_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 VDD a_1008_112# a_1028_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X15 a_960_156# a_544_476# a_644_576# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X16 VDD a_1008_112# a_2207_137# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 VSS TE a_36_137# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 VSS a_1008_112# a_2415_137# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X19 a_1008_112# a_644_576# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 VDD a_616_112# a_544_476# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_2415_137# CLK a_2207_137# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_2 CLK E Q TE VDD VSS
X0 VSS TE a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_975_112# a_682_576# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X2 a_682_576# a_582_476# a_462_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 VSS a_2159_122# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X4 a_314_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_2367_122# CLK a_2159_122# & Metric 1.00 nmos_6p0 w=1u l=0.6u
X6 a_682_576# a_572_112# a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X7 a_462_576# E a_314_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 VDD a_572_112# a_582_476# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X9 a_975_112# a_682_576# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 a_572_112# CLK VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 a_2159_122# CLK VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS a_975_112# a_916_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_984_576# a_572_112# a_682_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 VDD a_975_112# a_2159_122# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 Q a_2159_122# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X16 a_572_112# CLK VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 a_36_156# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 Q a_2159_122# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_916_156# a_582_476# a_682_576# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VDD a_2159_122# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VDD a_975_112# a_984_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 VSS a_572_112# a_582_476# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X23 VSS a_975_112# a_2367_122# & Metric 1.00 nmos_6p0 w=1u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__icgtp_4 CLK E Q TE VDD VSS
X0 VSS TE a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_572_112# CLK VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_964_112# a_692_156# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 VSS a_964_112# a_2356_133# & Metric 1.00 nmos_6p0 w=1u l=0.6u
X4 a_692_156# a_678_532# a_448_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_692_156# a_572_112# a_36_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 VSS a_2148_133# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X7 VDD a_572_112# a_678_532# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 a_964_112# a_692_156# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X9 a_2356_133# CLK a_2148_133# & Metric 1.00 nmos_6p0 w=1u l=0.6u
X10 a_572_112# CLK VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 VSS a_2148_133# Q & Metric 1.00 nmos_6p0 w=1u l=0.6u
X12 VSS a_572_112# a_678_532# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_984_576# a_572_112# a_692_156# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_2148_133# CLK VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VSS a_964_112# a_916_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X16 Q a_2148_133# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X17 a_36_156# E VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 VDD a_964_112# a_2148_133# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_300_576# TE VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 Q a_2148_133# VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X21 Q a_2148_133# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 Q a_2148_133# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_916_156# a_678_532# a_692_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 a_448_576# E a_300_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X25 VDD a_2148_133# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VDD a_2148_133# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD a_964_112# a_984_576# w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__icgtp_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_2 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_3 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_4 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_8 I VDD VSS ZN
X0 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_12 I VDD VSS ZN
X0 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_16 I VDD VSS ZN
X0 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_20.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_20 I VDD VSS ZN
X0 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 ZN I VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X35 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 ZN I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 VSS I ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 VDD I ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__inv_20.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_1 EN I VDD VSS ZN
X0 a_1368_171# I VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 a_517_215# a_36_215# a_428_683# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X2 VDD a_1368_171# a_428_683# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X3 VDD EN a_36_215# w_n86_453# pmos_6p0 w=0.99u l=0.5u
X4 a_428_683# EN a_517_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 VSS EN a_36_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 VDD a_428_683# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 a_428_683# EN VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X8 a_1368_171# I VDD w_n86_453# pmos_6p0 w=0.99u l=0.5u
X9 a_517_215# a_36_215# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 VSS a_1368_171# a_517_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X11 VSS a_517_215# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_2 EN I VDD VSS ZN
X0 a_951_24# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 VSS a_951_24# a_479_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_479_69# a_47_69# a_449_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VSS a_479_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_951_24# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_479_69# a_47_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN a_479_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD a_951_24# a_449_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X8 ZN a_449_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X9 VDD EN a_47_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 a_449_573# EN a_479_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD a_449_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 VSS EN a_47_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_449_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_3.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_3 EN I VDD VSS ZN
X0 ZN a_449_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 VSS I a_982_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN a_449_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VDD a_449_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X4 a_479_69# a_982_68# VSS & Metric 1.00 nmos_6p0 w=0.885u l=0.6u
X5 VDD I a_982_68# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 ZN a_479_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN a_479_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_479_69# a_47_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD EN a_47_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 a_449_573# a_982_68# VDD w_n86_453# pmos_6p0 w=1.485u l=0.5u
X11 a_449_573# EN a_479_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_479_69# a_47_69# a_449_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 VSS EN a_47_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 a_449_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 VSS a_982_68# a_479_69# & Metric 1.00 nmos_6p0 w=0.885u l=0.6u
X16 VSS a_479_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD a_982_68# a_449_573# w_n86_453# pmos_6p0 w=1.485u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_3.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_4 EN I VDD VSS ZN
X0 a_438_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 ZN a_438_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X2 ZN a_438_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VDD a_438_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X4 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD a_438_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VSS a_971_68# a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS I a_971_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_468_69# a_971_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_438_573# a_971_68# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X14 a_438_573# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD a_971_68# a_438_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X16 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD I a_971_68# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X18 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 a_468_69# a_36_69# a_438_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_8.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_8 EN I VDD VSS ZN
X0 a_556_573# a_1060_68# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD a_1060_68# a_556_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_468_68# a_1060_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_468_68# a_36_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_468_68# a_1060_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_556_573# EN a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VSS a_1060_68# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD a_556_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 VSS EN a_36_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 ZN a_556_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 VSS I a_1060_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 ZN a_556_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X17 VDD a_556_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X18 ZN a_556_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 VSS a_1060_68# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD a_556_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X21 a_556_573# a_1060_68# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X22 ZN a_556_573# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X23 VDD EN a_36_68# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X24 a_1060_68# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X25 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD a_556_573# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X27 a_556_573# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X28 VDD I a_1060_68# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X29 a_1060_68# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_468_68# a_36_68# a_556_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X32 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VDD a_1060_68# a_556_573# w_n86_453# pmos_6p0 w=1.8u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_8.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_12.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_12 EN I VDD VSS ZN
X0 a_468_69# a_36_69# a_541_575# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 VDD a_945_580# a_541_575# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X2 VSS a_945_580# a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS a_945_580# a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD a_945_580# a_541_575# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X7 a_468_69# a_945_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_541_575# a_945_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 a_541_575# a_945_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X12 a_945_580# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_468_69# a_945_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD a_945_580# a_541_575# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X16 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X17 a_468_69# a_945_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_541_575# a_945_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 a_468_69# a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_945_580# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X21 VSS I a_945_580# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 VSS I a_945_580# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 VDD I a_945_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X25 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X26 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X28 a_541_575# EN a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X30 VDD I a_945_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X31 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X32 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X33 VSS EN a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X35 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X36 VDD EN a_36_69# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X37 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X38 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 a_541_575# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X40 VDD a_541_575# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X41 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X42 VSS a_468_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VSS a_945_580# a_468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X44 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 ZN a_541_575# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X46 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X47 ZN a_468_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_12.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_16.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__invz_16 EN I VDD VSS ZN
X0 VDD I a_1108_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X1 a_468_68# a_1108_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_556_580# a_1108_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X3 VSS I a_1108_580# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X6 VSS I a_1108_580# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_468_68# a_36_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X10 VDD I a_1108_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X11 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X13 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X14 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X15 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X16 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 VDD a_1108_580# a_556_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X18 a_556_580# a_1108_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X19 a_556_580# EN a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD EN a_36_68# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X21 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X22 a_1108_580# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X23 VSS EN a_36_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VDD a_1108_580# a_556_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X26 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_556_580# EN VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X28 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 VDD a_1108_580# a_556_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X30 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_468_68# a_36_68# a_556_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X33 a_1108_580# I VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X34 a_556_580# a_1108_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X35 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X36 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X37 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X38 VSS a_1108_580# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 VSS a_1108_580# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 VSS a_1108_580# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X42 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X44 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 VDD a_1108_580# a_556_580# w_n86_453# pmos_6p0 w=1.8u l=0.5u
X46 a_468_68# a_1108_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X47 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X48 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X49 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X50 VSS a_1108_580# a_468_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X51 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
X52 a_1108_580# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X53 a_468_68# a_1108_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X54 VSS a_468_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X55 a_1108_580# I VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X56 ZN a_468_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X57 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X58 a_468_68# a_1108_580# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X59 a_556_580# a_1108_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X60 ZN a_556_580# VDD w_n86_453# pmos_6p0 w=1.8u l=0.5u
X61 VDD a_556_580# ZN w_n86_453# pmos_6p0 w=1.8u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__invz_16.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VSS
X0 a_1020_652# a_36_92# a_872_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_504_110# a_36_92# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_1364_532# a_1020_652# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 a_1224_652# a_504_110# a_1020_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 VSS a_1020_652# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_504_110# a_36_92# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD a_1020_652# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1264_107# a_36_92# a_1020_652# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 VSS E a_36_92# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 VSS a_1364_532# a_1264_107# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 VDD E a_36_92# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 VDD a_1364_532# a_1224_652# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_872_652# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_1364_532# a_1020_652# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_1020_652# a_504_110# a_872_107# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 a_872_107# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_2 D E Q VDD VSS
X0 a_1020_652# a_36_92# a_872_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_504_110# a_36_92# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 Q a_1020_652# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_1264_125# a_36_92# a_1020_652# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 a_1364_532# a_1020_652# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_1224_652# a_504_110# a_1020_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD a_1020_652# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 Q a_1020_652# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_504_110# a_36_92# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X9 VSS E a_36_92# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_1020_652# a_504_110# a_872_125# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 VSS a_1364_532# a_1264_125# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X12 VDD E a_36_92# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 VDD a_1364_532# a_1224_652# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_872_125# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 a_872_652# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VSS a_1020_652# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_1364_532# a_1020_652# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_4 D E Q VDD VSS
X0 VDD E a_37_134# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X1 Q a_1041_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS E a_37_134# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 VDD a_1041_69# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_933_649# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X5 VSS a_1041_69# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1041_69# a_37_134# a_933_649# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VSS a_1041_69# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_485_615# a_37_134# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_1265_69# a_37_134# a_1041_69# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 a_1285_649# a_485_615# a_1041_69# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_1405_25# a_1285_649# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 Q a_1041_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_1405_25# a_1041_69# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_1405_25# a_1041_69# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 Q a_1041_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD a_1041_69# a_1405_25# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 a_873_69# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 Q a_1041_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_1041_69# a_485_615# a_873_69# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 VSS a_1041_69# a_1405_25# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X21 VSS a_1405_25# a_1265_69# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_485_615# a_37_134# VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X23 VDD a_1041_69# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_1 D E Q RN VDD VSS
X0 a_672_157# D a_504_157# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X1 a_1112_113# a_388_674# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 VDD a_1112_113# a_1132_674# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_504_157# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 VDD E a_36_139# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_2018_598# a_1112_113# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 a_1232_157# a_1112_113# a_1064_157# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X7 VDD RN a_388_674# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 Q a_2018_598# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_780_674# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_1064_157# a_36_139# a_388_674# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 Q a_2018_598# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS E a_36_139# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X13 a_1112_113# a_388_674# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X14 a_388_674# a_36_139# a_780_674# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 a_388_674# E a_672_157# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X16 VSS RN a_1232_157# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 a_2018_598# a_1112_113# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_1132_674# E a_388_674# w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_2 D E Q RN VDD VSS
X0 VDD a_2059_598# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_409_736# a_61_138# a_801_736# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 a_2059_598# a_1153_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X3 a_1273_156# a_1153_112# a_1105_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 a_1153_736# E a_409_736# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_1105_156# a_61_138# a_409_736# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 VSS a_2059_598# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_545_156# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 a_2059_598# a_1153_112# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 a_1153_112# a_409_736# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 VDD a_1153_112# a_1153_736# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 Q a_2059_598# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD E a_61_138# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X13 VDD RN a_409_736# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_409_736# E a_713_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 VSS E a_61_138# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 a_713_156# D a_545_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 a_1153_112# a_409_736# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 Q a_2059_598# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS RN a_1273_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X20 a_801_736# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrnq_4 D E Q RN VDD VSS
X0 a_431_738# a_43_155# a_823_738# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VDD a_1195_112# a_2181_662# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X2 VDD a_2181_662# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_511_156# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 Q a_2181_662# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD E a_43_155# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X6 a_1239_738# E a_431_738# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VSS a_1195_112# a_2181_662# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 Q a_2181_662# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS RN a_1315_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 VSS a_431_738# a_1195_112# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X11 VSS a_2181_662# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD RN a_431_738# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_823_738# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_1315_156# a_1195_112# a_1147_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 VSS a_2181_662# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_2181_662# a_1195_112# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X17 a_1195_112# a_431_738# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X18 a_431_738# E a_679_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X19 VDD a_431_738# a_1195_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 VSS E a_43_155# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X21 a_2181_662# a_1195_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 Q a_2181_662# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_679_156# D a_511_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 a_1147_156# a_43_155# a_431_738# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X25 Q a_2181_662# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 VDD a_2181_662# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD a_1195_112# a_1239_738# w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_1195_112# a_431_738# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_1 D E Q RN SETN VDD VSS
X0 VDD RN a_396_648# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VDD a_1120_112# a_1140_648# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 a_680_156# D a_512_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X3 a_1668_156# a_396_648# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 VDD E a_36_138# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_788_648# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_1120_112# a_396_648# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_512_156# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 VSS E a_36_138# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 Q a_1996_175# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_1240_156# a_1120_112# a_1072_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X11 a_396_648# a_36_138# a_788_648# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_1072_156# a_36_138# a_396_648# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_1140_648# E a_396_648# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 VSS a_1120_112# a_1996_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 VDD SETN a_1120_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X16 a_396_648# E a_680_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X17 a_1120_112# SETN a_1668_156# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X18 Q a_1996_175# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VDD a_1120_112# a_1996_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 VSS RN a_1240_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_2 D E Q RN SETN VDD VSS
X0 a_1316_664# E a_404_740# w_n86_453# pmos_6p0 w=1u l=0.6u
X1 Q a_2128_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.6u
X2 VSS a_2128_69# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1324_156# a_1204_112# a_1156_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X4 VSS a_1204_112# a_2128_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD RN a_404_740# w_n86_453# pmos_6p0 w=1u l=0.6u
X6 a_404_740# a_36_664# a_924_664# w_n86_453# pmos_6p0 w=1u l=0.6u
X7 a_1156_156# a_36_664# a_404_740# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X8 VDD E a_36_664# w_n86_453# pmos_6p0 w=1.38u l=0.6u
X9 Q a_2128_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_1204_112# a_404_740# VDD w_n86_453# pmos_6p0 w=1u l=0.6u
X11 VDD a_1204_112# a_2128_69# w_n86_453# pmos_6p0 w=1.83u l=0.6u
X12 VDD SETN a_1204_112# w_n86_453# pmos_6p0 w=1.38u l=0.6u
X13 VSS E a_36_664# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 a_404_740# E a_764_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 a_1204_112# SETN a_1752_156# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 VDD a_2128_69# Q w_n86_453# pmos_6p0 w=1.83u l=0.6u
X17 a_548_156# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 VSS RN a_1324_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X19 a_924_664# D VDD w_n86_453# pmos_6p0 w=1u l=0.6u
X20 VDD a_1204_112# a_1316_664# w_n86_453# pmos_6p0 w=1u l=0.6u
X21 a_764_156# D a_548_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X22 a_1752_156# a_404_740# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latrsnq_4 D E Q RN SETN VDD VSS
X0 VDD a_1142_112# a_2216_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS RN a_1262_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 VSS a_2216_574# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1136_694# E a_392_694# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 VDD a_1142_112# a_1136_694# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 Q a_2216_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD a_2216_574# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS a_2216_574# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_1262_156# a_1142_112# a_1094_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X9 a_1142_112# a_392_694# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X10 VDD a_2216_574# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_1094_156# a_44_584# a_392_694# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X12 Q a_2216_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 Q a_2216_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_534_156# RN VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X15 a_2216_574# a_1142_112# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 VDD RN a_392_694# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 Q a_2216_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VSS E a_44_584# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 a_784_694# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X20 VDD E a_44_584# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 VSS a_1142_112# a_2216_574# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD SETN a_1142_112# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 a_392_694# E a_702_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 a_1142_112# SETN a_1690_156# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X25 a_392_694# a_44_584# a_784_694# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_702_156# D a_534_156# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X27 a_1690_156# a_392_694# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X28 a_2216_574# a_1142_112# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latrsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_1 D E Q SETN VDD VSS
X0 a_632_673# a_36_149# a_484_673# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VDD a_916_629# a_836_673# w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VSS a_916_629# a_896_167# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X3 a_836_673# E a_632_673# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_916_629# a_632_673# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_916_629# SETN a_1324_149# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 VSS a_916_629# a_1658_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 VDD SETN a_916_629# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 VSS E a_36_149# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 a_896_167# a_36_149# a_632_673# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X10 VDD a_916_629# a_1658_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X11 VDD E a_36_149# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_1324_149# a_632_673# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X13 a_632_673# E a_504_167# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X14 a_484_673# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X15 Q a_1658_175# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 Q a_1658_175# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_504_167# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_2 D E Q SETN VDD VSS
X0 a_894_653# a_642_697# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_894_653# a_896_134# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 VDD SETN a_894_653# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_494_697# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_896_134# a_36_134# a_642_697# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X5 Q a_1684_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD a_1684_69# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_1324_69# a_642_697# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_642_697# a_36_134# a_494_697# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 VSS a_894_653# a_1684_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VDD a_894_653# a_1684_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 a_894_653# SETN a_1324_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_642_697# E a_504_134# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X13 a_846_697# E a_642_697# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 Q a_1684_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD a_894_653# a_846_697# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VSS a_1684_69# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_504_134# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X18 VDD E a_36_134# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X19 VSS E a_36_134# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__latsnq_4 D E Q SETN VDD VSS
X0 a_533_708# D VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VSS a_949_664# a_911_192# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X2 a_1339_68# a_687_192# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_949_664# SETN a_1339_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_901_708# E a_687_192# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_911_192# a_51_174# a_687_192# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X6 VSS E a_51_174# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 VDD a_949_664# a_901_708# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 VSS a_949_664# a_1865_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 Q a_1865_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS a_1865_573# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_949_664# a_687_192# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1865_573# a_949_664# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS a_1865_573# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD a_1865_573# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD SETN a_949_664# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD a_949_664# a_1865_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 Q a_1865_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_687_192# E a_519_192# & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X19 VDD E a_51_174# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 a_1865_573# a_949_664# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD a_1865_573# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 Q a_1865_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_519_192# D VSS & Metric 1.00 nmos_6p0 w=0.7u l=0.6u
X24 Q a_1865_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_687_192# a_51_174# a_533_708# w_n86_453# pmos_6p0 w=1u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__latsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_1 I0 I1 S VDD VSS Z
X0 a_896_82# a_592_394# a_124_24# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 VSS I0 a_896_82# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 a_124_24# a_592_394# a_537_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_896_574# S a_124_24# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X4 a_504_82# I1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 a_124_24# S a_504_82# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 VSS a_124_24# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD I0 a_896_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X8 a_592_394# S VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X9 a_592_394# S VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X10 a_537_574# I1 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X11 VDD a_124_24# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_2 I0 I1 S VDD VSS Z
X0 a_848_529# S VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_124_25# a_848_529# a_692_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS I0 a_1084_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1152_573# S a_124_25# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_1084_69# a_848_529# a_124_25# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS a_124_25# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_692_69# I1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD a_124_25# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD I0 a_1152_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_124_25# S a_692_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_124_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_692_573# I1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_848_529# S VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 Z a_124_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux2_4 I0 I1 S VDD VSS Z
X0 a_1307_529# S VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VDD a_135_25# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_135_25# S a_1151_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1151_573# I1 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_1543_69# a_1307_529# a_135_25# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD a_135_25# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_135_25# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VSS a_135_25# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_1151_69# I1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_135_25# a_1307_529# a_1151_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_1611_573# S a_135_25# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 Z a_135_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 Z a_135_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VSS I0 a_1543_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD I0 a_1611_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 Z a_135_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1307_529# S VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 Z a_135_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_1 I0 I1 I2 I3 S0 S1 VDD VSS Z
X0 a_234_669# I2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 Z a_1056_112# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X2 a_692_156# S0 a_468_156# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X3 a_2362_201# I1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 VSS I0 a_2770_669# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 a_1056_112# S1 a_468_156# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 VDD S1 a_1436_481# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X7 a_2362_201# I1 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X8 a_2770_669# a_348_112# a_1740_669# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X9 a_1056_112# a_1436_481# a_468_156# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X10 a_1740_669# a_348_112# a_2362_201# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X11 a_2770_669# S0 a_1740_669# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X12 a_348_112# S0 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X13 a_1740_669# S1 a_1056_112# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X14 a_468_156# a_348_112# a_234_669# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X15 a_348_112# S0 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X16 VSS S1 a_1436_481# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X17 VDD I0 a_2770_669# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X18 VDD I3 a_692_156# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X19 VSS I3 a_692_156# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X20 a_468_156# S0 a_234_669# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X21 a_1740_669# a_1436_481# a_1056_112# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X22 a_1740_669# S0 a_2362_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X23 a_692_156# a_348_112# a_468_156# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X24 a_234_669# I2 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X25 Z a_1056_112# VSS & Metric 1.00 nmos_6p0 w=0.9u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_2 I0 I1 I2 I3 S0 S1 VDD VSS Z
X0 a_758_596# a_484_112# a_516_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X1 a_1156_112# a_1861_464# a_516_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X2 a_244_156# I2 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X3 a_244_156# I2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X4 a_2195_156# a_1861_464# a_1156_112# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X5 a_3209_596# a_484_112# a_2195_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X6 VDD I0 a_3209_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X7 a_484_112# S0 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X8 VSS a_1156_112# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X9 VSS S1 a_1861_464# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 a_516_596# S0 a_244_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X11 a_758_596# S0 a_516_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X12 a_2195_156# S0 a_2787_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X13 a_2195_156# S1 a_1156_112# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X14 a_3209_596# S0 a_2195_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X15 a_516_596# a_484_112# a_244_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X16 VSS I0 a_3209_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 Z a_1156_112# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X18 VDD S1 a_1861_464# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X19 a_2195_156# a_484_112# a_2787_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X20 a_1156_112# S1 a_516_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X21 Z a_1156_112# VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X22 a_484_112# S0 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X23 VDD a_1156_112# Z w_n86_453# pmos_6p0 w=1.28u l=0.5u
X24 a_2787_156# I1 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X25 a_2787_156# I1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X26 VDD I3 a_758_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X27 VSS I3 a_758_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__mux4_4 I0 I1 I2 I3 S0 S1 VDD VSS Z
X0 a_2596_156# a_2360_496# a_1169_115# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X1 VDD a_1169_115# Z w_n86_453# pmos_6p0 w=1.28u l=0.5u
X2 a_1169_115# a_2360_496# a_529_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X3 a_497_115# S0 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X4 Z a_1169_115# VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X5 a_2596_156# S1 a_1169_115# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X6 a_3236_156# I1 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X7 VDD a_1169_115# Z w_n86_453# pmos_6p0 w=1.28u l=0.5u
X8 a_3236_156# I1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X9 a_257_159# I2 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X10 VSS I3 a_755_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X11 a_257_159# I2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X12 VDD S1 a_2360_496# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X13 VDD I3 a_755_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X14 a_3684_156# a_497_115# a_2596_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X15 Z a_1169_115# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X16 a_1169_115# S1 a_529_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X17 a_3684_156# S0 a_2596_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X18 a_755_596# a_497_115# a_529_596# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X19 VDD I0 a_3684_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X20 VSS a_1169_115# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X21 a_529_596# S0 a_257_159# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X22 a_497_115# S0 VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X23 VSS S1 a_2360_496# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X24 a_755_596# S0 a_529_596# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X25 a_2596_156# S0 a_3236_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X26 a_2596_156# a_497_115# a_3236_156# w_n86_453# pmos_6p0 w=1.28u l=0.5u
X27 a_529_596# a_497_115# a_257_159# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X28 Z a_1169_115# VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X29 Z a_1169_115# VSS & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X30 VSS a_1169_115# Z & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
X31 VSS I0 a_3684_156# & Metric 1.00 nmos_6p0 w=0.8u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__mux4_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_1 A1 A2 VDD VSS ZN
X0 ZN A2 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X1 VDD A1 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X2 ZN A1 a_245_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_245_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_2 A1 A2 VDD VSS ZN
X0 a_652_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS A2 a_652_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A2 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X3 VDD A1 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X4 ZN A1 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X5 VDD A2 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X6 ZN A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand2_4 A1 A2 VDD VSS ZN
X0 ZN A1 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN A2 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X2 a_661_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_1060_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD A1 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X5 a_260_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN A1 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X7 VSS A2 a_1468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD A2 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X9 ZN A2 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X10 VSS A2 a_661_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD A1 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X12 ZN A1 a_260_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_1468_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 ZN A1 VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X15 VDD A2 ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_1 A1 A2 A3 VDD VSS ZN
X0 ZN A3 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 VDD A2 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 a_271_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_455_69# A2 a_271_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN A1 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X5 ZN A1 a_455_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_2 A1 A2 A3 VDD VSS ZN
X0 a_856_68# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VDD A1 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 a_272_68# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN A2 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X4 VDD A3 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X5 ZN A1 a_448_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_1040_68# A2 a_856_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN A3 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X8 a_448_68# A2 a_272_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS A3 a_1040_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VDD A2 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X11 ZN A1 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand3_4 A1 A2 A3 VDD VSS ZN
X0 VDD A1 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 ZN A1 a_1732_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A2 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X3 VSS A3 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS A3 a_1100_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD A3 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X6 VDD A1 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X7 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_672_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN A2 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X10 ZN A3 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X11 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD A2 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X13 ZN A1 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X14 VDD A3 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X15 a_36_69# A2 a_672_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 ZN A1 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X17 a_1732_69# A2 a_1528_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_244_69# A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 ZN A3 VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X20 a_1528_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD A2 ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X22 a_1100_69# A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand3_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_1 A1 A2 A3 A4 VDD VSS ZN
X0 VDD A3 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X1 ZN A2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X2 VDD A1 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X3 a_275_69# A4 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_673_69# A2 a_469_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_469_69# A3 a_275_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN A1 a_673_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN A4 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_2 A1 A2 A3 A4 VDD VSS ZN
X0 ZN A1 a_632_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN A2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X2 VDD A3 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X3 a_1060_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_1254_69# A2 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN A4 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X6 VSS A4 a_1458_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD A4 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X8 a_1458_69# A3 a_1254_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN A3 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X10 a_632_69# A2 a_438_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD A2 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X12 a_244_69# A4 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 ZN A1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X14 VDD A1 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X15 a_438_69# A3 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nand4_4 A1 A2 A3 A4 VDD VSS ZN
X0 a_652_69# A4 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_36_69# A3 a_652_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD A4 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X3 VSS A4 a_1060_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN A4 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X5 a_1060_69# A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_36_69# A2 a_3100_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD A3 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X8 ZN A1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X9 ZN A2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X10 VDD A2 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X11 VDD A1 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X12 a_36_69# A2 a_2284_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 ZN A3 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X14 a_1662_69# A3 a_1468_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_2284_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 ZN A2 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X17 ZN A1 a_1866_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD A2 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X19 VDD A4 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X20 VDD A1 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X21 ZN A4 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X22 ZN A1 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X23 VSS A4 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_2692_69# A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 ZN A1 a_2692_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 a_244_69# A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_1468_69# A4 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 VDD A3 ZN w_n86_453# pmos_6p0 w=1.28u l=0.5u
X29 a_1866_69# A2 a_1662_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 ZN A3 VDD w_n86_453# pmos_6p0 w=1.28u l=0.5u
X31 a_3100_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nand4_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_1 A1 A2 VDD VSS ZN
X0 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X1 ZN A1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X3 a_234_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_2 A1 A2 VDD VSS ZN
X0 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X1 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X2 a_672_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X4 ZN A1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X6 a_234_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VDD A2 a_672_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor2_4 A1 A2 VDD VSS ZN
X0 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X1 a_682_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X3 ZN A1 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X5 ZN A1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X7 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X8 a_1130_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VDD A2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X11 a_1578_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X13 a_234_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.92u l=0.6u
X15 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_1 A1 A2 A3 VDD VSS ZN
X0 ZN A1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_244_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_2 A1 A2 A3 VDD VSS ZN
X0 ZN A1 a_468_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_468_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 VDD A3 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 a_1130_573# A2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_244_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X11 a_906_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor3_4 A1 A2 A3 VDD VSS ZN
X0 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X1 a_1568_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_224_573# A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_672_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 ZN A1 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 VDD A3 a_1120_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN A1 a_1792_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X12 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X13 a_1792_573# A2 a_1568_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X15 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X16 VDD A3 a_224_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 a_1120_573# A2 a_36_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X21 a_36_573# A2 a_672_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 a_36_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor3_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_1 A1 A2 A3 A4 VDD VSS ZN
X0 a_682_573# A2 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X3 a_458_573# A3 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_244_573# A4 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 ZN A4 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X7 ZN A1 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_2 A1 A2 A3 A4 VDD VSS ZN
X0 ZN A1 a_1213_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_683_573# A4 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X3 a_1213_573# A2 a_943_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 a_943_573# A3 a_683_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS A4 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X7 a_1661_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X9 a_57_573# A2 a_1661_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN A4 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X11 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X12 VDD A4 a_245_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X14 a_245_573# A3 a_57_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__nor4_4 A1 A2 A3 A4 VDD VSS ZN
X0 VDD A4 a_1265_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X3 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_3793_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_745_573# A4 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_3273_573# A2 a_119_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS A4 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X8 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X9 a_1265_573# A3 a_119_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_119_573# A3 a_745_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 ZN A1 a_2233_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 ZN A1 a_3273_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS A1 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X14 ZN A4 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X15 VSS A2 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X16 a_2233_573# A2 a_1973_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_2753_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X19 ZN A4 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X20 a_1973_573# A3 a_1713_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_119_573# A2 a_2753_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_119_573# A2 a_3793_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VDD A4 a_307_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 ZN A3 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X25 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X26 a_1713_573# A4 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VSS A3 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X28 ZN A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X29 a_307_573# A3 a_119_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 ZN A1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X31 VSS A4 ZN & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__nor4_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_1 A1 A2 B VDD VSS ZN
X0 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X2 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN A1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_234_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_2 A1 A2 B VDD VSS ZN
X0 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X1 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X3 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD A2 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_1130_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_692_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 ZN A1 a_692_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai21_4 A1 A2 B VDD VSS ZN
X0 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_682_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN A1 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN A1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X7 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X8 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X11 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_1130_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VDD A2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_244_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X17 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_1578_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai21_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_1 A1 A2 B1 B2 VDD VSS ZN
X0 a_682_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN B1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_244_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_2 A1 A2 B1 B2 VDD VSS ZN
X0 a_682_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A1 a_1140_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_1140_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD A2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_244_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN B1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_1578_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD B2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai22_4 A1 A2 B1 B2 VDD VSS ZN
X0 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_2474_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VDD A2 a_3370_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 ZN B1 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_3370_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN A1 a_2036_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_1130_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_2922_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD B2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD A2 a_2474_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 ZN B1 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 a_1578_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_692_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 a_234_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 ZN A1 a_2922_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 VDD B2 a_692_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_2036_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai22_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_1 A1 A2 A3 B VDD VSS ZN
X0 a_682_573# A2 a_468_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_468_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN A3 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X5 a_244_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_244_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD A3 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_2 A1 A2 A3 B VDD VSS ZN
X0 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_1354_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X4 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X5 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 ZN A1 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VDD A3 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1578_573# A2 a_1354_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_692_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_906_573# A2 a_692_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai31_4 A1 A2 A3 B VDD VSS ZN
X0 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X1 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD A3 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_2474_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN A1 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_2026_573# A2 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X9 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_56_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VDD B ZN w_n86_453# pmos_6p0 w=1.645u l=0.5u
X12 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_56_573# A2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN B VDD w_n86_453# pmos_6p0 w=1.645u l=0.5u
X15 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_36_69# B VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 ZN A1 a_2026_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 a_1130_573# A2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 VDD A3 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VSS B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 a_1578_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_906_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_56_573# A2 a_2474_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai31_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_1 A1 A2 A3 B1 B2 VDD VSS ZN
X0 ZN A1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VSS A2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_244_69# B2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_244_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_244_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_244_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD B2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_906_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_2 A1 A2 A3 B1 B2 VDD VSS ZN
X0 ZN A1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_36_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_2026_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_36_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_36_69# B2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_36_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD A3 a_1120_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_36_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_1588_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 ZN B1 a_1588_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_244_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD B2 a_2026_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VSS A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1120_573# A2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 ZN B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 ZN B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_906_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai32_4 A1 A2 A3 B1 B2 VDD VSS ZN
X0 a_77_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN A1 a_87_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_275_573# A2 a_87_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_87_573# A2 a_733_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_77_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_77_69# B2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_77_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_77_69# B2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_1619_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS A2 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN B2 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_733_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_77_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_3515_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN B2 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VSS A3 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_77_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 ZN B1 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_87_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 ZN B1 a_3077_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 VSS A2 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 ZN B1 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_3963_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VDD B2 a_4411_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VSS A1 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VSS A3 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD A3 a_1171_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 ZN A1 a_1843_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_4411_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 VSS A1 a_77_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 a_77_69# B1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_1171_573# A2 a_87_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X32 a_1843_573# A2 a_1619_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 a_77_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 ZN B1 a_3963_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 a_3077_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 a_77_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 VDD A3 a_275_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X38 VDD B2 a_3515_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 a_87_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai32_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_1 A1 A2 A3 B1 B2 B3 VDD VSS ZN
X0 ZN B1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 ZN A3 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD A3 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_458_573# B2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_244_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_1130_573# A2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_244_573# B3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_244_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_244_69# B3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_906_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_2 A1 A2 A3 B1 B2 B3 VDD VSS ZN
X0 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN B1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_2474_573# A2 a_2250_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD B3 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN A1 a_1802_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_36_69# B3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_458_573# B2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_1588_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_2250_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_1130_573# B2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_1802_573# A2 a_1588_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_244_573# B3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS B3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_906_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VDD A3 a_2474_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai33_4 A1 A2 A3 B1 B2 B3 VDD VSS ZN
X0 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_2848_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_682_573# B3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN B1 a_1802_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_36_69# B3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD A3 a_4818_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_3922_573# A2 a_3698_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_36_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD B3 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_2848_573# A2 a_5266_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_3698_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_36_69# B3 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_1130_573# B2 a_46_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_36_69# A3 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 a_1802_573# B2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_5266_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 VDD A3 a_3922_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_4818_573# A2 a_2848_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 ZN A1 a_2848_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 VSS B3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 VDD B3 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 a_1578_573# B3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 a_46_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X37 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 a_2848_573# A2 a_4380_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 VSS B1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 ZN A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 ZN B1 a_46_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X42 ZN A1 a_2848_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X43 a_234_573# B2 a_46_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X44 VSS B3 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 a_46_573# B2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X46 a_46_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X47 a_4380_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai33_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_1 A1 A2 B C VDD VSS ZN
X0 VDD B ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 VSS C a_698_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_698_69# B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_244_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_2 A1 A2 B C VDD VSS ZN
X0 VSS C a_1146_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_682_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_1146_69# B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 ZN A1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_244_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN B VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X8 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X9 a_1564_69# C VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_36_69# B a_1564_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X14 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD B ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai211_4 A1 A2 B C VDD VSS ZN
X0 VSS C a_2868_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_682_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X3 a_2042_69# B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X5 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN A1 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN B VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X8 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN A1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VDD B ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X11 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X12 ZN B VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X13 VDD B ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X14 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X16 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 a_2868_69# B a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_36_69# B a_3276_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_1130_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VSS C a_2042_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 VDD A2 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_244_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 a_1578_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_36_69# B a_2460_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 a_2460_69# C VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X30 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_3276_69# C VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai211_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_1 A1 A2 B1 B2 C VDD VSS ZN
X0 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 a_36_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 ZN A2 a_698_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_698_69# C a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_244_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_698_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 ZN B1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_928_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS B2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN A1 a_928_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_2 A1 A2 B1 B2 C VDD VSS ZN
X0 a_36_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X2 ZN A2 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_474_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_2044_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 ZN A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN B1 a_474_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_244_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_36_69# C a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_36_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD A2 a_1606_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_244_69# C a_36_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VSS B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X16 VDD B2 a_912_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 a_1606_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN A1 a_2044_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_912_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai221_4 A1 A2 B1 B2 C VDD VSS ZN
X0 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X1 a_682_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_1972_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VDD B2 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_1972_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 ZN A1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VDD A2 a_3076_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_3962_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_244_69# C a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1972_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 ZN A1 a_4410_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN A1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 ZN A2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VSS B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_4410_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD B2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_244_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 ZN A2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VDD C ZN w_n86_453# pmos_6p0 w=1.46u l=0.5u
X22 a_1972_69# C a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_1130_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X25 ZN B1 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_244_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X27 VDD A2 a_3962_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X28 a_1972_69# C a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X29 a_3076_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 ZN A1 a_3524_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_1972_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 a_1578_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 a_244_69# B1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X35 a_3524_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 ZN C VDD w_n86_453# pmos_6p0 w=1.46u l=0.5u
X37 a_244_69# B2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X38 ZN B1 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 a_244_69# C a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai221_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_1 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 a_244_69# B1 a_628_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 a_628_69# B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VSS C1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN C1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VDD B2 a_826_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_628_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_244_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_826_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_1284_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_244_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN A1 a_1284_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 ZN A2 a_628_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_2 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 ZN B1 a_1722_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_682_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 ZN A2 a_1076_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_2170_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 ZN A1 a_2618_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_1722_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS C1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_1076_69# B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS C2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD C2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_1076_69# B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1076_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD B2 a_1274_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_244_573# C1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_1076_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_244_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_244_69# B2 a_1076_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_2618_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_244_69# C1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_244_69# B1 a_1076_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 VDD A2 a_2170_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 ZN C1 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 ZN A1 a_1076_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_1274_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__oai222_4 A1 A2 B1 B2 C1 C2 VDD VSS ZN
X0 a_682_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_2180_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_1972_69# B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN A2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_3514_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_1972_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS C1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD C2 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_1972_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD A2 a_4858_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS C2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_244_69# B1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD B2 a_3066_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_3962_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_244_69# B2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_1972_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_1972_69# A1 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 ZN A1 a_4410_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 ZN B1 a_2618_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 ZN A1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_244_69# B2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VSS C1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_4410_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 VSS C2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X24 VDD C2 a_234_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 a_244_69# C1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 ZN A2 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_1972_69# B1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 a_1130_573# C1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 ZN C1 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 VDD A2 a_3962_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X31 a_1972_69# B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_4858_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 ZN A1 a_5306_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X34 ZN B1 a_3514_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 a_244_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X36 a_1972_69# B2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 a_1578_573# C2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X38 a_2618_573# B2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X39 a_244_69# C1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X40 a_5306_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X41 a_234_573# C1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X42 VDD B2 a_2180_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X43 a_244_69# C2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X44 ZN A1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X45 ZN C1 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X46 a_3066_573# B1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X47 a_244_69# B1 a_1972_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__oai222_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1 A1 A2 VDD VSS Z
X0 a_255_756# A1 a_67_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 VSS A2 a_67_756# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X2 VDD A2 a_255_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 Z a_67_756# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_67_756# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_67_756# A1 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_2 A1 A2 VDD VSS Z
X0 Z a_56_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_56_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VSS A2 a_56_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_244_573# A1 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 Z a_56_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_56_573# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD a_56_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_4 A1 A2 VDD VSS Z
X0 a_682_573# A1 a_244_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A2 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VSS A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_244_69# A1 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_244_573# A2 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_244_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD A2 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or3_1 A1 A2 A3 VDD VSS Z
X0 Z a_36_101# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS A3 a_36_101# & Metric 1.00 nmos_6p0 w=0.525u l=0.6u
X2 a_36_101# A2 VSS & Metric 1.00 nmos_6p0 w=0.525u l=0.6u
X3 a_458_756# A2 a_244_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X4 a_244_756# A1 a_36_101# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X5 Z a_36_101# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS A1 a_36_101# & Metric 1.00 nmos_6p0 w=0.525u l=0.6u
X7 VDD A3 a_458_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or3_2 A1 A2 A3 VDD VSS Z
X0 VDD A3 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VDD a_36_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 Z a_36_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_36_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_36_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X5 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_244_573# A1 a_36_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS A3 a_36_69# & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X8 VSS A1 a_36_69# & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X9 VSS a_36_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or3_4 A1 A2 A3 VDD VSS Z
X0 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 a_244_69# A1 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS A3 a_244_69# & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X4 VSS A1 a_244_69# & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X5 VDD A3 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VSS A2 a_244_69# & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X9 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X11 a_1130_573# A2 a_906_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_244_573# A3 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 a_244_69# A1 VSS & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X16 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_244_69# A3 VSS & Metric 1.00 nmos_6p0 w=1.05u l=0.6u
X18 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_906_573# A1 a_244_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or3_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or4_1 A1 A2 A3 A4 VDD VSS Z
X0 a_484_756# A2 a_244_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 VSS A2 a_56_756# & Metric 1.00 nmos_6p0 w=0.395u l=0.6u
X2 a_718_756# A3 a_484_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_244_756# A1 a_56_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X4 VDD A4 a_718_756# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X5 VSS A4 a_56_756# & Metric 1.00 nmos_6p0 w=0.395u l=0.6u
X6 a_56_756# A1 VSS & Metric 1.00 nmos_6p0 w=0.395u l=0.6u
X7 Z a_56_756# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_56_756# A3 VSS & Metric 1.00 nmos_6p0 w=0.395u l=0.6u
X9 Z a_56_756# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or4_2 A1 A2 A3 A4 VDD VSS Z
X0 a_682_573# A3 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS a_56_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 VSS A4 a_56_573# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 VSS A2 a_56_573# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X4 a_458_573# A2 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_244_573# A1 a_56_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD a_56_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_56_573# A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X8 a_56_573# A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X9 Z a_56_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 Z a_56_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VDD A4 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__or4_4 A1 A2 A3 A4 VDD VSS Z
X0 a_682_573# A2 a_458_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS A4 a_244_69# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X2 a_1354_573# A2 a_1130_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS A2 a_244_69# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 VSS A1 a_244_69# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X6 VSS A3 a_244_69# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 a_458_573# A3 a_244_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_244_69# A1 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1130_573# A1 a_244_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 VDD A4 a_1578_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_244_573# A4 VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 VSS a_244_69# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X16 a_244_69# A2 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X17 a_1578_573# A3 a_1354_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 a_244_69# A4 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X19 VDD a_244_69# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 Z a_244_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 Z a_244_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 a_244_69# A3 VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 a_244_69# A1 a_682_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__or4_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_1 CLK D Q SE SI VDD VSS
X0 a_1712_582# a_1193_582# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X1 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 a_3276_608# a_3014_652# VSS & Metric 1.00 nmos_6p0 w=0.75u l=0.6u
X3 a_2332_226# a_1712_582# a_2098_652# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X4 a_800_652# SE a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_445_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD D a_800_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_2380_182# a_2098_652# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X8 VSS a_3276_608# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X10 a_3228_652# a_1712_582# a_3014_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_3276_608# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_2098_652# a_1193_582# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X13 VSS a_3276_608# a_3248_226# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X14 VDD a_3276_608# a_3228_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 a_2312_652# a_1193_582# a_2098_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_3014_652# a_1712_582# a_2380_182# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X17 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X18 VSS a_2380_182# a_2332_226# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X19 VSS CLK a_1193_582# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_2380_182# a_2098_652# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X21 a_2098_652# a_1712_582# a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 a_3276_608# a_3014_652# VDD w_n86_453# pmos_6p0 w=1.1u l=0.5u
X23 a_596_652# a_36_156# a_445_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_3014_652# a_1193_582# a_2380_182# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 VSS D a_860_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X26 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 VDD a_2380_182# a_2312_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_1712_582# a_1193_582# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X29 a_3248_226# a_1193_582# a_3014_652# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X30 VDD CLK a_1193_582# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X31 a_860_156# a_36_156# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_2 CLK D Q SE SI VDD VSS
X0 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X1 VSS a_2392_172# a_2344_216# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 VSS a_3400_24# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD a_3400_24# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_2392_172# a_2120_216# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X5 VSS a_3400_24# a_3260_216# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_468_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_626_652# a_36_156# a_468_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_3260_216# a_1232_174# a_3026_652# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X9 a_2120_216# a_1752_174# a_626_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_2470_652# a_1232_174# a_2120_216# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 Q a_3400_24# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X13 VSS CLK a_1232_174# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 a_2344_216# a_1752_174# a_2120_216# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X15 a_3240_652# a_1752_174# a_3026_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 VDD CLK a_1232_174# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X19 a_1752_174# a_1232_174# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X20 VDD a_3400_24# a_3240_652# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 VDD D a_850_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X22 a_1752_174# a_1232_174# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 VDD a_2392_172# a_2470_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_3400_24# a_3026_652# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X25 Q a_3400_24# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_2392_172# a_2120_216# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 VSS D a_860_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X28 a_850_652# SE a_626_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 a_2120_216# a_1232_174# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X30 a_3400_24# a_3026_652# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_3026_652# a_1232_174# a_2392_172# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_860_156# a_36_156# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X33 a_3026_652# a_1752_174# a_2392_172# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffq_4 CLK D Q SE SI VDD VSS
X0 Q a_3400_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X2 a_1752_175# a_1232_175# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X3 a_2440_652# a_1232_175# a_2120_217# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_2120_217# a_1232_175# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X5 a_3400_25# a_3026_652# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_3400_25# a_3026_652# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 VDD a_2392_173# a_2440_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_2392_173# a_2120_217# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_3026_652# a_1752_175# a_2392_173# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X10 VSS a_2392_173# a_2344_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X11 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X12 a_2392_173# a_2120_217# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X13 Q a_3400_25# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_3240_652# a_1752_175# a_3026_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 VDD CLK a_1232_175# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X16 a_2120_217# a_1752_175# a_652_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 VSS a_3400_25# a_3260_217# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VDD a_3400_25# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X20 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X21 a_1752_175# a_1232_175# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_3260_217# a_1232_175# a_3026_652# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X23 VDD a_3400_25# a_3240_652# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X24 VSS a_3400_25# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VDD D a_856_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_504_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 VSS a_3400_25# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X28 a_652_652# a_36_156# a_504_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 VDD a_3400_25# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X30 Q a_3400_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 VSS D a_860_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X32 VSS CLK a_1232_175# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X33 a_2344_217# a_1752_175# a_2120_217# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X34 a_856_652# SE a_652_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X35 a_3026_652# a_1232_175# a_2392_173# w_n86_453# pmos_6p0 w=1u l=0.5u
X36 Q a_3400_25# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 a_860_156# a_36_156# a_636_156# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1 CLK D Q RN SE SI VDD VSS
X0 a_468_187# SI VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X1 VSS a_3491_141# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_3116_185# a_1220_166# a_2292_141# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_840_652# D a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_2412_185# a_2292_141# a_2244_185# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X5 VSS a_3491_141# a_3340_185# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X6 a_1632_589# a_1220_166# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 a_3340_185# a_1632_589# a_3116_185# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_2292_141# a_1994_652# VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X9 VDD SE a_840_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_2198_652# a_1220_166# a_1994_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_2292_141# a_1994_652# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_1994_652# a_1220_166# a_636_187# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X13 VDD a_3491_141# a_3340_185# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 VSS a_36_187# a_860_187# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X15 a_1994_652# a_1632_589# a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_3340_185# a_1220_166# a_3116_185# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X17 VDD CLK a_1220_166# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X18 a_3491_141# a_3116_185# a_3835_185# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X19 a_3491_141# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X20 a_860_187# D a_636_187# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X21 VSS SE a_36_187# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X22 VSS CLK a_1220_166# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X23 VDD a_3116_185# a_3491_141# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 VDD a_2292_141# a_2198_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_2244_185# a_1632_589# a_1994_652# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X26 a_2198_652# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_448_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_3116_185# a_1632_589# a_2292_141# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X29 a_596_652# a_36_187# a_448_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_636_187# SE a_468_187# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X31 VDD SE a_36_187# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 VDD a_3491_141# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 VSS RN a_2412_185# & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
X34 a_1632_589# a_1220_166# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X35 a_3835_185# RN VSS & Metric 1.00 nmos_6p0 w=0.58u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2 CLK D Q RN SE SI VDD VSS
X0 a_2173_652# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 Q a_3421_151# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_3045_195# a_1621_580# a_2277_608# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_840_652# D a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_3273_195# a_1229_166# a_3045_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 VDD CLK a_1229_166# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 a_3421_151# a_3045_195# a_3801_124# & Metric 1.00 nmos_6p0 w=1u l=0.6u
X8 VDD SE a_840_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 a_1621_580# a_1229_166# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X10 a_1969_652# a_1229_166# a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X11 a_3801_124# RN VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X12 a_2425_195# a_2277_608# a_2257_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 a_2277_608# a_1969_652# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 a_3421_151# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X16 a_1621_580# a_1229_166# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X17 a_2257_195# a_1621_580# a_1969_652# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_3045_195# a_1229_166# a_2277_608# w_n86_453# pmos_6p0 w=1u l=0.5u
X20 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 VSS a_3421_151# a_3273_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 VDD a_3045_195# a_3421_151# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X23 VSS RN a_2425_195# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_3273_195# a_1621_580# a_3045_195# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_448_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X26 Q a_3421_151# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_2277_608# a_1969_652# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_596_652# a_36_156# a_448_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 VDD a_3421_151# a_3273_195# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_2173_652# a_1229_166# a_1969_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X31 VSS a_36_156# a_860_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X32 VDD a_3421_151# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X33 VDD a_2277_608# a_2173_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X34 a_1969_652# a_1621_580# a_596_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X35 a_860_156# D a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X36 VSS CLK a_1229_166# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X37 VSS a_3421_151# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4 CLK D Q RN SE SI VDD VSS
X0 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 a_724_156# SE a_556_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 a_2332_652# a_1312_163# a_2128_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_2128_652# a_1312_163# a_724_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_3432_206# a_1312_163# a_3208_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X5 a_3540_162# a_3208_206# a_3920_124# & Metric 1.00 nmos_6p0 w=1u l=0.6u
X6 VDD a_2436_608# a_2332_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VSS a_36_156# a_948_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_556_156# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_1714_580# a_1312_163# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X10 a_2332_652# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_3208_206# a_1312_163# a_2436_608# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_536_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X13 VDD a_3540_162# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_3208_206# a_1714_580# a_2436_608# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 VSS RN a_2592_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 VSS a_3540_162# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X17 a_684_652# a_36_156# a_536_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 VDD a_3540_162# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS a_3540_162# a_3432_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X20 Q a_3540_162# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 a_2436_608# a_2128_652# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X22 Q a_3540_162# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_2592_206# a_2436_608# a_2424_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_3920_124# RN VSS & Metric 1.00 nmos_6p0 w=1u l=0.6u
X25 VDD CLK a_1312_163# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 a_948_156# D a_724_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_3432_206# a_1714_580# a_3208_206# w_n86_453# pmos_6p0 w=1u l=0.5u
X28 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 VSS CLK a_1312_163# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X30 a_1714_580# a_1312_163# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X31 a_928_652# D a_684_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 VSS a_3540_162# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X33 VDD a_3540_162# a_3432_206# w_n86_453# pmos_6p0 w=1u l=0.5u
X34 VDD a_3208_206# a_3540_162# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X35 Q a_3540_162# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 Q a_3540_162# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X37 VDD SE a_928_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X38 a_3540_162# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X39 a_2436_608# a_2128_652# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X40 a_2128_652# a_1714_580# a_684_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X41 a_2424_206# a_1714_580# a_2128_652# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1 CLK D Q RN SE SETN SI VDD VSS
X0 VSS a_41_157# a_865_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 a_3600_215# a_1200_584# a_3376_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 a_4008_157# SETN a_3600_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 VDD a_3376_215# a_4056_113# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X4 a_1592_584# a_1200_584# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_3600_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD CLK a_1200_584# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X7 a_4400_157# RN VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 a_865_157# D a_641_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_1592_584# a_1200_584# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X10 a_2148_591# a_1200_584# a_1944_591# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VSS SE a_41_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X12 VDD a_2252_547# a_2148_591# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_4056_113# a_3376_215# a_4400_157# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X14 VSS RN a_2432_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 a_2984_215# a_1944_591# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 a_1944_591# a_1592_584# a_591_651# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 VDD SE a_41_157# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_3376_215# a_1592_584# a_2252_547# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 a_443_651# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X20 a_2252_547# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X21 VSS CLK a_1200_584# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X22 a_591_651# a_41_157# a_443_651# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 a_3376_215# a_1200_584# a_2252_547# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_1944_591# a_1200_584# a_641_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_641_157# SE a_473_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X26 VSS a_4056_113# a_4008_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_2148_591# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 VDD a_1944_591# a_2252_547# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 a_845_651# D a_591_651# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 Q a_4056_113# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_3600_215# a_1592_584# a_3376_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 VDD SE a_845_651# w_n86_453# pmos_6p0 w=1u l=0.5u
X33 a_2432_215# a_2252_547# a_2264_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X34 a_473_157# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X35 Q a_4056_113# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X36 a_2252_547# SETN a_2984_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X37 a_2264_215# a_1592_584# a_1944_591# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X38 VDD a_4056_113# a_3600_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X39 a_4056_113# RN VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2 CLK D Q RN SE SETN SI VDD VSS
X0 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 a_1972_588# a_1232_608# a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 VDD a_1972_588# a_2280_544# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_4008_157# SETN a_3600_226# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 VSS CLK a_1232_608# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_2948_226# a_1972_588# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 a_3600_226# a_1232_608# a_3376_226# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X7 a_840_652# D a_606_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X8 a_2480_226# a_2280_544# a_2312_226# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_4400_157# RN VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 VSS a_4056_113# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VDD SE a_840_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 a_2176_588# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X13 a_2280_544# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_2312_226# a_1624_608# a_1972_588# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_3376_226# a_1232_608# a_2280_544# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 VDD a_4056_113# a_3600_226# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 a_458_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X20 VDD CLK a_1232_608# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X21 a_3376_226# a_1624_608# a_2280_544# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_3600_226# a_1624_608# a_3376_226# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VSS RN a_2480_226# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_3600_226# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_1624_608# a_1232_608# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X26 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 VSS a_4056_113# a_4008_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 VDD a_3376_226# a_4056_113# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X29 a_1624_608# a_1232_608# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X30 Q a_4056_113# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X31 a_4056_113# a_3376_226# a_4400_157# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_606_652# a_36_156# a_458_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X33 a_2176_588# a_1232_608# a_1972_588# w_n86_453# pmos_6p0 w=1u l=0.5u
X34 VDD a_4056_113# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X35 VSS a_36_156# a_860_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X36 VDD a_2280_544# a_2176_588# w_n86_453# pmos_6p0 w=1u l=0.5u
X37 a_4056_113# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X38 a_1972_588# a_1624_608# a_606_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X39 Q a_4056_113# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X40 a_2280_544# SETN a_2948_226# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X41 a_860_156# D a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4 CLK D Q RN SE SETN SI VDD VSS
X0 a_2931_215# a_1955_577# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 VDD a_3323_215# a_4049_137# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD SE a_36_199# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_2463_215# a_2263_533# a_2295_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_3323_215# a_1127_596# a_2263_533# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_636_199# SE a_468_199# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 a_428_652# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_3323_215# a_1607_596# a_2263_533# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 VDD a_4049_137# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_576_652# a_36_199# a_428_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X10 a_3547_215# a_1607_596# a_3323_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X11 a_2295_215# a_1607_596# a_1955_577# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X12 a_4049_137# RN VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 Q a_4049_137# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_780_652# D a_576_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 a_468_199# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X16 Q a_4049_137# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS a_4049_137# a_4001_181# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X18 a_4049_137# a_3323_215# a_4393_181# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_1607_596# a_1127_596# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 VDD a_4049_137# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_1607_596# a_1127_596# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X22 a_2159_577# RN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X23 VSS RN a_2463_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 Q a_4049_137# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VDD a_4049_137# a_3547_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 VSS a_36_199# a_860_199# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_2263_533# SETN a_2931_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 VDD SE a_780_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X29 a_860_199# D a_636_199# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X30 VDD CLK a_1127_596# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X31 a_2159_577# a_1127_596# a_1955_577# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_3547_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X33 VSS SE a_36_199# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X34 a_3547_215# a_1127_596# a_3323_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X35 a_4001_181# SETN a_3547_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X36 VSS a_4049_137# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X37 VDD a_2263_533# a_2159_577# w_n86_453# pmos_6p0 w=1u l=0.5u
X38 a_2263_533# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X39 VSS CLK a_1127_596# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X40 VSS a_4049_137# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X41 a_1955_577# a_1607_596# a_576_652# w_n86_453# pmos_6p0 w=1u l=0.5u
X42 Q a_4049_137# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X43 VDD a_1955_577# a_2263_533# w_n86_453# pmos_6p0 w=1u l=0.5u
X44 a_1955_577# a_1127_596# a_636_199# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X45 a_4393_181# RN VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffrsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1 CLK D Q SE SETN SI VDD VSS
X0 a_3430_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X1 VSS a_36_206# a_860_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 a_840_644# D a_596_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X3 a_3430_215# a_1274_158# a_3206_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X4 a_2064_582# a_1686_577# a_596_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X5 a_860_206# D a_636_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X6 a_3994_160# a_3206_215# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X7 a_1686_577# a_1274_158# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X8 VSS SE a_36_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X9 a_2064_582# a_1274_158# a_636_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X10 a_3206_215# a_1686_577# a_2346_113# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X11 VDD CLK a_1274_158# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X12 a_1686_577# a_1274_158# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X13 a_3946_204# SETN a_3430_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X14 VSS a_2346_113# a_2298_157# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 VDD SE a_840_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X16 a_3994_160# a_3206_215# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X17 VDD a_2346_113# a_2278_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 a_636_206# SE a_468_206# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X19 a_2298_157# a_1686_577# a_2064_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X20 a_448_644# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X21 Q a_3994_160# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X22 Q a_3994_160# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_596_644# a_36_206# a_448_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X24 a_2278_582# a_1274_158# a_2064_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X25 a_3206_215# a_1274_158# a_2346_113# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 VSS CLK a_1274_158# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X27 a_2346_113# a_2064_582# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_468_206# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 VDD SE a_36_206# w_n86_453# pmos_6p0 w=1u l=0.5u
X30 VDD SETN a_2346_113# w_n86_453# pmos_6p0 w=1u l=0.5u
X31 a_3430_215# a_1686_577# a_3206_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 VDD a_3994_160# a_3430_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X33 a_2778_215# a_2064_582# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X34 a_2346_113# SETN a_2778_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X35 VSS a_3994_160# a_3946_204# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2 CLK D Q SE SETN SI VDD VSS
X0 a_2239_582# a_1235_164# a_2025_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X1 a_3327_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X2 VSS a_2307_130# a_2259_174# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X3 VDD SE a_855_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X4 a_1647_573# a_1235_164# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X5 a_2307_130# a_2025_582# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X6 VDD a_3927_171# a_3327_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X7 a_2695_215# a_2025_582# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X8 VDD SETN a_2307_130# w_n86_453# pmos_6p0 w=1u l=0.5u
X9 Q a_3927_171# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 Q a_3927_171# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 VSS a_51_196# a_875_196# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X12 a_2259_174# a_1647_573# a_2025_582# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X13 a_3927_171# a_3103_215# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD SE a_51_196# w_n86_453# pmos_6p0 w=1u l=0.5u
X15 a_3927_171# a_3103_215# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD a_2307_130# a_2239_582# w_n86_453# pmos_6p0 w=1u l=0.5u
X17 a_3327_215# a_1647_573# a_3103_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X18 VDD a_3927_171# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X19 VSS CLK a_1235_164# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X20 a_3103_215# a_1647_573# a_2307_130# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X21 VSS a_3927_171# a_3863_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_2025_582# a_1647_573# a_641_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X23 a_875_196# D a_651_196# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 VSS SE a_51_196# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_3103_215# a_1235_164# a_2307_130# w_n86_453# pmos_6p0 w=1u l=0.5u
X26 a_3863_215# SETN a_3327_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X27 a_855_644# D a_641_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X28 a_2307_130# SETN a_2695_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_483_644# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X30 a_651_196# SE a_483_196# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X31 a_641_644# a_51_196# a_483_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X32 a_2025_582# a_1235_164# a_651_196# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X33 VSS a_3927_171# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X34 a_1647_573# a_1235_164# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X35 a_3327_215# a_1235_164# a_3103_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X36 VDD CLK a_1235_164# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X37 a_483_196# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4 CLK D Q SE SETN SI VDD VSS
X0 VSS SE a_36_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X1 a_2236_476# SETN a_2684_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X2 a_3861_140# a_3076_215# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS a_3076_215# a_3861_140# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS CLK a_1224_166# & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X5 a_840_644# D a_596_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X6 a_3300_215# SETN VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X7 VDD a_3076_215# a_3861_140# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 VDD a_3861_140# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 VSS a_3861_140# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_445_644# SI VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X11 VDD a_2236_476# a_2188_577# w_n86_453# pmos_6p0 w=1u l=0.5u
X12 VDD SE a_840_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X13 VDD a_3861_140# a_3300_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X14 a_2684_215# a_1984_577# VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X15 Q a_3861_140# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_2236_476# a_1984_577# VDD w_n86_453# pmos_6p0 w=1u l=0.5u
X17 VDD a_3861_140# Q w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VDD SETN a_2236_476# w_n86_453# pmos_6p0 w=1u l=0.5u
X19 Q a_3861_140# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X20 a_3861_140# a_3076_215# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X21 VSS a_3861_140# a_3813_184# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X22 a_636_156# SE a_468_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X23 VSS a_2236_476# a_2248_154# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X24 a_1984_577# a_1224_166# a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X25 a_3813_184# SETN a_3300_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X26 a_3076_215# a_1224_166# a_2236_476# w_n86_453# pmos_6p0 w=1u l=0.5u
X27 a_468_156# SI VSS & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X28 a_3076_215# a_1626_608# a_2236_476# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X29 a_1626_608# a_1224_166# VSS & Metric 1.00 nmos_6p0 w=0.79u l=0.6u
X30 a_3300_215# a_1626_608# a_3076_215# w_n86_453# pmos_6p0 w=1u l=0.5u
X31 Q a_3861_140# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X32 a_596_644# a_36_156# a_445_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X33 VDD CLK a_1224_166# w_n86_453# pmos_6p0 w=1.38u l=0.5u
X34 VSS a_36_156# a_860_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X35 VDD SE a_36_156# w_n86_453# pmos_6p0 w=1u l=0.5u
X36 a_2188_577# a_1224_166# a_1984_577# w_n86_453# pmos_6p0 w=1u l=0.5u
X37 a_2248_154# a_1626_608# a_1984_577# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X38 Q a_3861_140# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X39 a_1626_608# a_1224_166# VDD w_n86_453# pmos_6p0 w=1.38u l=0.5u
X40 a_3300_215# a_1224_166# a_3076_215# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X41 a_1984_577# a_1626_608# a_596_644# w_n86_453# pmos_6p0 w=1u l=0.5u
X42 a_860_156# D a_636_156# & Metric 1.00 nmos_6p0 w=0.59u l=0.6u
X43 VSS a_3861_140# Q & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__sdffsnq_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__tieh.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__tieh VDD VSS Z
X0 Z a_125_157# VDD w_n86_453# pmos_6p0 w=0.9u l=0.5u
X1 a_125_157# a_125_157# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__tieh.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__tiel.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__tiel VDD VSS ZN
X0 ZN a_124_157# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 a_124_157# a_124_157# VDD w_n86_453# pmos_6p0 w=0.9u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__tiel.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_1 A1 A2 VDD VSS ZN
X0 a_44_201# A2 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 VDD A1 a_44_201# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X2 a_696_69# A2 ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 VDD A2 a_910_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS A1 a_252_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X5 a_696_69# a_44_201# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_910_573# A1 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 ZN a_44_201# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 ZN A1 a_696_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_252_201# A2 a_44_201# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_2 A1 A2 VDD VSS ZN
X0 a_728_69# a_56_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 ZN a_728_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VSS A2 a_952_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 a_952_69# A1 a_728_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS a_728_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS A1 a_56_574# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 ZN a_728_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_728_574# a_56_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X8 a_728_69# A1 a_728_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_56_574# A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X10 VDD A1 a_244_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X11 a_244_574# A2 a_56_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X12 a_728_574# A2 a_728_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 VDD a_728_69# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor2_4 A1 A2 VDD VSS ZN
X0 a_728_69# a_46_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X1 VSS A2 a_952_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_952_69# A1 a_728_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X3 ZN a_728_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 VSS a_728_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_728_69# A1 a_708_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 VDD A1 a_234_573# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X7 VSS A1 a_46_573# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 VSS a_728_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 ZN a_728_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 a_708_573# A2 a_728_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 ZN a_728_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD a_728_69# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 ZN a_728_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 a_708_573# a_46_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD a_728_69# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_234_573# A2 a_46_573# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X17 a_46_573# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_1 A1 A2 A3 VDD VSS ZN
X0 a_244_691# A2 a_56_691# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X1 a_718_691# a_56_691# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X2 a_718_691# A2 a_728_146# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_728_146# a_56_691# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_1296_146# a_728_146# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X5 a_1948_69# a_1296_146# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD A3 a_1296_146# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X7 a_1504_146# a_728_146# a_1296_146# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X8 a_56_691# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 VSS A2 a_952_146# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X10 a_1948_69# a_728_146# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 ZN a_1296_146# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_952_146# A1 a_728_146# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X13 a_2172_573# A3 ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X14 ZN A3 a_1948_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X15 VDD a_728_146# a_2172_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_728_146# A1 a_718_691# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X17 VSS A3 a_1504_146# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X18 VDD A1 a_244_691# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X19 VSS A1 a_56_691# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_2 A1 A2 A3 VDD VSS ZN
X0 a_752_702# A2 a_752_167# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 VDD A3 a_1528_704# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X2 a_2002_573# a_1340_704# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS A3 a_1340_704# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_268_705# A2 a_80_705# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X5 VSS a_2012_68# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VSS A2 a_976_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X7 a_80_705# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 a_2236_68# A3 a_2012_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_2012_68# a_1340_704# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X10 ZN a_2012_68# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_1340_704# a_752_167# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X12 a_976_167# A1 a_752_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X13 VDD A1 a_268_705# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X14 a_2012_68# A3 a_2002_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 a_2002_573# a_752_167# a_2012_68# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 a_752_702# a_80_705# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X17 ZN a_2012_68# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 VSS a_752_167# a_2236_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 VSS A1 a_80_705# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X20 a_752_167# A1 a_752_702# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X21 a_752_167# a_80_705# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X22 a_1528_704# a_752_167# a_1340_704# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X23 VDD a_2012_68# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xnor3_4 A1 A2 A3 VDD VSS ZN
X0 a_1307_678# a_692_167# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X1 a_56_705# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X2 a_1987_573# a_692_167# a_1987_69# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS a_1987_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 a_1987_573# a_1307_678# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 ZN a_1987_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_692_678# a_56_705# VDD w_n86_453# pmos_6p0 w=0.495u l=0.5u
X7 a_692_167# a_56_705# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X8 a_692_167# A1 a_692_678# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X9 VDD a_1987_69# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 VSS A2 a_916_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X11 a_1495_678# a_692_167# a_1307_678# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X12 VSS a_692_167# a_2211_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_2211_69# A3 a_1987_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VDD A3 a_1495_678# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X15 ZN a_1987_69# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VSS A3 a_1307_678# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X17 VSS A1 a_56_705# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X18 ZN a_1987_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_692_678# A2 a_692_167# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X20 VDD a_1987_69# ZN w_n86_453# pmos_6p0 w=1.83u l=0.5u
X21 a_916_167# A1 a_692_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X22 ZN a_1987_69# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X23 a_244_705# A2 a_56_705# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X24 a_1987_69# a_1307_678# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X25 VSS a_1987_69# ZN & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X26 VDD A1 a_244_705# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X27 a_1987_69# A3 a_1987_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xnor3_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_1 A1 A2 VDD VSS Z
X0 VSS A1 a_56_573# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X1 Z A1 a_718_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 VDD A1 a_244_573# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_244_573# A2 a_56_573# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X4 a_718_573# a_56_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_718_573# A2 Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X6 a_56_573# A2 VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X7 Z a_56_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 VSS A2 a_952_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_952_68# A1 Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_2 A1 A2 VDD VSS Z
X0 VDD A1 a_36_166# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X1 a_688_69# A2 a_678_574# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X2 a_912_574# A1 a_678_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VSS A1 a_244_166# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X4 a_688_69# a_36_166# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 VSS a_678_574# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 VDD A2 a_912_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_678_574# A1 a_688_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X8 Z a_678_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 a_244_166# A2 a_36_166# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X10 a_678_574# a_36_166# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 Z a_678_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X12 a_36_166# A2 VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X13 VDD a_678_574# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor2_4 A1 A2 VDD VSS Z
X0 a_688_573# a_36_260# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X1 VDD A2 a_902_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 a_902_573# A1 a_688_573# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_688_573# A1 a_688_68# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 Z a_688_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X5 a_244_260# A2 a_36_260# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X6 VSS a_688_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X7 a_36_260# A2 VDD w_n86_453# pmos_6p0 w=0.495u l=0.5u
X8 VSS a_688_573# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X9 VDD A1 a_36_260# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X10 Z a_688_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 Z a_688_573# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD a_688_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X13 a_688_68# A2 a_688_573# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 Z a_688_573# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X15 VDD a_688_573# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VSS A1 a_244_260# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X17 a_688_68# a_36_260# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor2_4.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_1.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_1 A1 A2 A3 VDD VSS Z
X0 VDD A1 a_244_642# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X1 VSS A1 a_56_642# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X2 VDD A3 a_1501_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X3 a_2212_69# A3 Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X4 VSS a_728_166# a_2212_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_728_166# a_56_642# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 Z A3 a_1978_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 VSS A3 a_1313_574# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X8 a_1978_574# a_728_166# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X9 a_1501_574# a_728_166# a_1313_574# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X10 a_1313_574# a_728_166# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X11 a_56_642# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X12 VSS A2 a_952_166# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X13 a_728_166# A1 a_718_642# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X14 a_244_642# A2 a_56_642# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X15 a_718_642# a_56_642# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X16 a_718_642# A2 a_728_166# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X17 a_1978_574# a_1313_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X18 Z a_1313_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_952_166# A1 a_728_166# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_1.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_2.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_2 A1 A2 A3 VDD VSS Z
X0 VDD A1 a_244_700# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X1 a_728_167# A1 a_718_616# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X2 a_2172_574# A3 a_1938_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 VDD a_1938_574# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X4 a_56_700# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X5 VSS A2 a_952_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X6 VDD a_728_167# a_2172_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X7 a_244_700# A2 a_56_700# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X8 a_718_616# a_56_700# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X9 a_718_616# A2 a_728_167# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X10 a_1948_69# a_1296_167# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X11 a_952_167# A1 a_728_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X12 a_1948_69# a_728_167# a_1938_574# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X13 a_1296_167# a_728_167# VDD w_n86_453# pmos_6p0 w=0.915u l=0.5u
X14 VDD A3 a_1296_167# w_n86_453# pmos_6p0 w=0.915u l=0.5u
X15 Z a_1938_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VSS A3 a_1504_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X17 Z a_1938_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X18 VSS A1 a_56_700# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X19 a_1938_574# A3 a_1948_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X20 a_728_167# a_56_700# VSS & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
X21 VSS a_1938_574# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X22 a_1938_574# a_1296_167# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X23 a_1504_167# a_728_167# a_1296_167# & Metric 1.00 nmos_6p0 w=0.66u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_2.ext - technology: gf180mcuC



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_4.ext - technology: gf180mcuC

.subckt gf180mcu_fd_sc_mcu9t5v0__xor3_4 A1 A2 A3 VDD VSS Z
X0 a_692_710# a_56_737# VDD w_n86_453# pmos_6p0 w=0.495u l=0.5u
X1 a_2126_574# A3 a_1912_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X2 Z a_1912_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X3 a_56_737# A2 VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X4 VSS a_1912_574# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X5 a_1912_69# a_692_167# a_1912_574# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X6 a_692_167# A1 a_692_710# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X7 a_1260_167# a_692_167# VDD w_n86_453# pmos_6p0 w=0.495u l=0.5u
X8 a_692_167# a_56_737# VSS & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X9 VDD a_1912_574# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X10 Z a_1912_574# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X11 VSS a_1912_574# Z & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X12 VDD A3 a_1260_167# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X13 Z a_1912_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X14 VSS A3 a_1468_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X15 a_1912_574# a_1260_167# VDD w_n86_453# pmos_6p0 w=1.83u l=0.5u
X16 VDD a_1912_574# Z w_n86_453# pmos_6p0 w=1.83u l=0.5u
X17 VSS A2 a_916_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X18 Z a_1912_574# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X19 a_692_710# A2 a_692_167# w_n86_453# pmos_6p0 w=0.495u l=0.5u
X20 a_244_737# A2 a_56_737# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X21 VSS A1 a_56_737# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X22 VDD A1 a_244_737# w_n86_453# pmos_6p0 w=0.36u l=0.5u
X23 a_1468_167# a_692_167# a_1260_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X24 a_916_167# A1 a_692_167# & Metric 1.00 nmos_6p0 w=0.36u l=0.6u
X25 VDD a_692_167# a_2126_574# w_n86_453# pmos_6p0 w=1.83u l=0.5u
X26 a_1912_574# A3 a_1912_69# & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
X27 a_1912_69# a_1260_167# VSS & Metric 1.00 nmos_6p0 w=1.32u l=0.6u
.ends



******* EOF

* NGSPICE file created from gf180mcu_fd_sc_mcu9t5v0__xor3_4.ext - technology: gf180mcuC



******* EOF

