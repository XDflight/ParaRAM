magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 2170 27755 10792 29293
<< mvnmos >>
rect 4129 26006 4269 27006
rect 5191 26006 5331 27006
rect 5435 26006 5575 27006
rect 5679 26006 5819 27006
rect 5923 26006 6063 27006
rect 6167 26006 6307 27006
rect 6411 26006 6551 27006
rect 6655 26006 6795 27006
rect 6899 26006 7039 27006
rect 7143 26006 7283 27006
rect 7387 26006 7527 27006
rect 7631 26006 7771 27006
rect 7875 26006 8015 27006
<< mvpmos >>
rect 2665 27917 2805 28917
rect 2909 27917 3049 28917
rect 3153 27917 3293 28917
rect 3397 27917 3537 28917
rect 3641 27917 3781 28917
rect 3885 27917 4025 28917
rect 4129 27917 4269 28917
rect 4545 27917 4685 28917
rect 4789 27917 4929 28917
rect 5033 27917 5173 28917
rect 5277 27917 5417 28917
rect 5521 27917 5661 28917
rect 5765 27917 5905 28917
rect 6009 27917 6149 28917
rect 6253 27917 6393 28917
rect 6497 27917 6637 28917
rect 6741 27917 6881 28917
rect 6985 27917 7125 28917
rect 7229 27917 7369 28917
rect 7473 27917 7613 28917
rect 7717 27917 7857 28917
rect 7961 27917 8101 28917
rect 8205 27917 8345 28917
rect 8449 27917 8589 28917
rect 8693 27917 8833 28917
rect 8937 27917 9077 28917
rect 9181 27917 9321 28917
rect 9425 27917 9565 28917
rect 9669 27917 9809 28917
rect 9913 27917 10053 28917
rect 10157 27917 10297 28917
<< mvndiff >>
rect 4041 26993 4129 27006
rect 4041 26947 4054 26993
rect 4100 26947 4129 26993
rect 4041 26890 4129 26947
rect 4041 26844 4054 26890
rect 4100 26844 4129 26890
rect 4041 26787 4129 26844
rect 4041 26741 4054 26787
rect 4100 26741 4129 26787
rect 4041 26684 4129 26741
rect 4041 26638 4054 26684
rect 4100 26638 4129 26684
rect 4041 26581 4129 26638
rect 4041 26535 4054 26581
rect 4100 26535 4129 26581
rect 4041 26478 4129 26535
rect 4041 26432 4054 26478
rect 4100 26432 4129 26478
rect 4041 26375 4129 26432
rect 4041 26329 4054 26375
rect 4100 26329 4129 26375
rect 4041 26272 4129 26329
rect 4041 26226 4054 26272
rect 4100 26226 4129 26272
rect 4041 26169 4129 26226
rect 4041 26123 4054 26169
rect 4100 26123 4129 26169
rect 4041 26065 4129 26123
rect 4041 26019 4054 26065
rect 4100 26019 4129 26065
rect 4041 26006 4129 26019
rect 4269 26993 4357 27006
rect 4269 26947 4298 26993
rect 4344 26947 4357 26993
rect 4269 26890 4357 26947
rect 4269 26844 4298 26890
rect 4344 26844 4357 26890
rect 4269 26787 4357 26844
rect 4269 26741 4298 26787
rect 4344 26741 4357 26787
rect 4269 26684 4357 26741
rect 4269 26638 4298 26684
rect 4344 26638 4357 26684
rect 4269 26581 4357 26638
rect 4269 26535 4298 26581
rect 4344 26535 4357 26581
rect 4269 26478 4357 26535
rect 4269 26432 4298 26478
rect 4344 26432 4357 26478
rect 4269 26375 4357 26432
rect 4269 26329 4298 26375
rect 4344 26329 4357 26375
rect 4269 26272 4357 26329
rect 4269 26226 4298 26272
rect 4344 26226 4357 26272
rect 4269 26169 4357 26226
rect 4269 26123 4298 26169
rect 4344 26123 4357 26169
rect 4269 26065 4357 26123
rect 4269 26019 4298 26065
rect 4344 26019 4357 26065
rect 4269 26006 4357 26019
rect 5103 26993 5191 27006
rect 5103 26947 5116 26993
rect 5162 26947 5191 26993
rect 5103 26890 5191 26947
rect 5103 26844 5116 26890
rect 5162 26844 5191 26890
rect 5103 26787 5191 26844
rect 5103 26741 5116 26787
rect 5162 26741 5191 26787
rect 5103 26684 5191 26741
rect 5103 26638 5116 26684
rect 5162 26638 5191 26684
rect 5103 26581 5191 26638
rect 5103 26535 5116 26581
rect 5162 26535 5191 26581
rect 5103 26478 5191 26535
rect 5103 26432 5116 26478
rect 5162 26432 5191 26478
rect 5103 26375 5191 26432
rect 5103 26329 5116 26375
rect 5162 26329 5191 26375
rect 5103 26272 5191 26329
rect 5103 26226 5116 26272
rect 5162 26226 5191 26272
rect 5103 26169 5191 26226
rect 5103 26123 5116 26169
rect 5162 26123 5191 26169
rect 5103 26065 5191 26123
rect 5103 26019 5116 26065
rect 5162 26019 5191 26065
rect 5103 26006 5191 26019
rect 5331 26993 5435 27006
rect 5331 26947 5360 26993
rect 5406 26947 5435 26993
rect 5331 26890 5435 26947
rect 5331 26844 5360 26890
rect 5406 26844 5435 26890
rect 5331 26787 5435 26844
rect 5331 26741 5360 26787
rect 5406 26741 5435 26787
rect 5331 26684 5435 26741
rect 5331 26638 5360 26684
rect 5406 26638 5435 26684
rect 5331 26581 5435 26638
rect 5331 26535 5360 26581
rect 5406 26535 5435 26581
rect 5331 26478 5435 26535
rect 5331 26432 5360 26478
rect 5406 26432 5435 26478
rect 5331 26375 5435 26432
rect 5331 26329 5360 26375
rect 5406 26329 5435 26375
rect 5331 26272 5435 26329
rect 5331 26226 5360 26272
rect 5406 26226 5435 26272
rect 5331 26169 5435 26226
rect 5331 26123 5360 26169
rect 5406 26123 5435 26169
rect 5331 26065 5435 26123
rect 5331 26019 5360 26065
rect 5406 26019 5435 26065
rect 5331 26006 5435 26019
rect 5575 26993 5679 27006
rect 5575 26947 5604 26993
rect 5650 26947 5679 26993
rect 5575 26890 5679 26947
rect 5575 26844 5604 26890
rect 5650 26844 5679 26890
rect 5575 26787 5679 26844
rect 5575 26741 5604 26787
rect 5650 26741 5679 26787
rect 5575 26684 5679 26741
rect 5575 26638 5604 26684
rect 5650 26638 5679 26684
rect 5575 26581 5679 26638
rect 5575 26535 5604 26581
rect 5650 26535 5679 26581
rect 5575 26478 5679 26535
rect 5575 26432 5604 26478
rect 5650 26432 5679 26478
rect 5575 26375 5679 26432
rect 5575 26329 5604 26375
rect 5650 26329 5679 26375
rect 5575 26272 5679 26329
rect 5575 26226 5604 26272
rect 5650 26226 5679 26272
rect 5575 26169 5679 26226
rect 5575 26123 5604 26169
rect 5650 26123 5679 26169
rect 5575 26065 5679 26123
rect 5575 26019 5604 26065
rect 5650 26019 5679 26065
rect 5575 26006 5679 26019
rect 5819 26993 5923 27006
rect 5819 26947 5848 26993
rect 5894 26947 5923 26993
rect 5819 26890 5923 26947
rect 5819 26844 5848 26890
rect 5894 26844 5923 26890
rect 5819 26787 5923 26844
rect 5819 26741 5848 26787
rect 5894 26741 5923 26787
rect 5819 26684 5923 26741
rect 5819 26638 5848 26684
rect 5894 26638 5923 26684
rect 5819 26581 5923 26638
rect 5819 26535 5848 26581
rect 5894 26535 5923 26581
rect 5819 26478 5923 26535
rect 5819 26432 5848 26478
rect 5894 26432 5923 26478
rect 5819 26375 5923 26432
rect 5819 26329 5848 26375
rect 5894 26329 5923 26375
rect 5819 26272 5923 26329
rect 5819 26226 5848 26272
rect 5894 26226 5923 26272
rect 5819 26169 5923 26226
rect 5819 26123 5848 26169
rect 5894 26123 5923 26169
rect 5819 26065 5923 26123
rect 5819 26019 5848 26065
rect 5894 26019 5923 26065
rect 5819 26006 5923 26019
rect 6063 26993 6167 27006
rect 6063 26947 6092 26993
rect 6138 26947 6167 26993
rect 6063 26890 6167 26947
rect 6063 26844 6092 26890
rect 6138 26844 6167 26890
rect 6063 26787 6167 26844
rect 6063 26741 6092 26787
rect 6138 26741 6167 26787
rect 6063 26684 6167 26741
rect 6063 26638 6092 26684
rect 6138 26638 6167 26684
rect 6063 26581 6167 26638
rect 6063 26535 6092 26581
rect 6138 26535 6167 26581
rect 6063 26478 6167 26535
rect 6063 26432 6092 26478
rect 6138 26432 6167 26478
rect 6063 26375 6167 26432
rect 6063 26329 6092 26375
rect 6138 26329 6167 26375
rect 6063 26272 6167 26329
rect 6063 26226 6092 26272
rect 6138 26226 6167 26272
rect 6063 26169 6167 26226
rect 6063 26123 6092 26169
rect 6138 26123 6167 26169
rect 6063 26065 6167 26123
rect 6063 26019 6092 26065
rect 6138 26019 6167 26065
rect 6063 26006 6167 26019
rect 6307 26993 6411 27006
rect 6307 26947 6336 26993
rect 6382 26947 6411 26993
rect 6307 26890 6411 26947
rect 6307 26844 6336 26890
rect 6382 26844 6411 26890
rect 6307 26787 6411 26844
rect 6307 26741 6336 26787
rect 6382 26741 6411 26787
rect 6307 26684 6411 26741
rect 6307 26638 6336 26684
rect 6382 26638 6411 26684
rect 6307 26581 6411 26638
rect 6307 26535 6336 26581
rect 6382 26535 6411 26581
rect 6307 26478 6411 26535
rect 6307 26432 6336 26478
rect 6382 26432 6411 26478
rect 6307 26375 6411 26432
rect 6307 26329 6336 26375
rect 6382 26329 6411 26375
rect 6307 26272 6411 26329
rect 6307 26226 6336 26272
rect 6382 26226 6411 26272
rect 6307 26169 6411 26226
rect 6307 26123 6336 26169
rect 6382 26123 6411 26169
rect 6307 26065 6411 26123
rect 6307 26019 6336 26065
rect 6382 26019 6411 26065
rect 6307 26006 6411 26019
rect 6551 26993 6655 27006
rect 6551 26947 6580 26993
rect 6626 26947 6655 26993
rect 6551 26890 6655 26947
rect 6551 26844 6580 26890
rect 6626 26844 6655 26890
rect 6551 26787 6655 26844
rect 6551 26741 6580 26787
rect 6626 26741 6655 26787
rect 6551 26684 6655 26741
rect 6551 26638 6580 26684
rect 6626 26638 6655 26684
rect 6551 26581 6655 26638
rect 6551 26535 6580 26581
rect 6626 26535 6655 26581
rect 6551 26478 6655 26535
rect 6551 26432 6580 26478
rect 6626 26432 6655 26478
rect 6551 26375 6655 26432
rect 6551 26329 6580 26375
rect 6626 26329 6655 26375
rect 6551 26272 6655 26329
rect 6551 26226 6580 26272
rect 6626 26226 6655 26272
rect 6551 26169 6655 26226
rect 6551 26123 6580 26169
rect 6626 26123 6655 26169
rect 6551 26065 6655 26123
rect 6551 26019 6580 26065
rect 6626 26019 6655 26065
rect 6551 26006 6655 26019
rect 6795 26993 6899 27006
rect 6795 26947 6824 26993
rect 6870 26947 6899 26993
rect 6795 26890 6899 26947
rect 6795 26844 6824 26890
rect 6870 26844 6899 26890
rect 6795 26787 6899 26844
rect 6795 26741 6824 26787
rect 6870 26741 6899 26787
rect 6795 26684 6899 26741
rect 6795 26638 6824 26684
rect 6870 26638 6899 26684
rect 6795 26581 6899 26638
rect 6795 26535 6824 26581
rect 6870 26535 6899 26581
rect 6795 26478 6899 26535
rect 6795 26432 6824 26478
rect 6870 26432 6899 26478
rect 6795 26375 6899 26432
rect 6795 26329 6824 26375
rect 6870 26329 6899 26375
rect 6795 26272 6899 26329
rect 6795 26226 6824 26272
rect 6870 26226 6899 26272
rect 6795 26169 6899 26226
rect 6795 26123 6824 26169
rect 6870 26123 6899 26169
rect 6795 26065 6899 26123
rect 6795 26019 6824 26065
rect 6870 26019 6899 26065
rect 6795 26006 6899 26019
rect 7039 26993 7143 27006
rect 7039 26947 7068 26993
rect 7114 26947 7143 26993
rect 7039 26890 7143 26947
rect 7039 26844 7068 26890
rect 7114 26844 7143 26890
rect 7039 26787 7143 26844
rect 7039 26741 7068 26787
rect 7114 26741 7143 26787
rect 7039 26684 7143 26741
rect 7039 26638 7068 26684
rect 7114 26638 7143 26684
rect 7039 26581 7143 26638
rect 7039 26535 7068 26581
rect 7114 26535 7143 26581
rect 7039 26478 7143 26535
rect 7039 26432 7068 26478
rect 7114 26432 7143 26478
rect 7039 26375 7143 26432
rect 7039 26329 7068 26375
rect 7114 26329 7143 26375
rect 7039 26272 7143 26329
rect 7039 26226 7068 26272
rect 7114 26226 7143 26272
rect 7039 26169 7143 26226
rect 7039 26123 7068 26169
rect 7114 26123 7143 26169
rect 7039 26065 7143 26123
rect 7039 26019 7068 26065
rect 7114 26019 7143 26065
rect 7039 26006 7143 26019
rect 7283 26993 7387 27006
rect 7283 26947 7312 26993
rect 7358 26947 7387 26993
rect 7283 26890 7387 26947
rect 7283 26844 7312 26890
rect 7358 26844 7387 26890
rect 7283 26787 7387 26844
rect 7283 26741 7312 26787
rect 7358 26741 7387 26787
rect 7283 26684 7387 26741
rect 7283 26638 7312 26684
rect 7358 26638 7387 26684
rect 7283 26581 7387 26638
rect 7283 26535 7312 26581
rect 7358 26535 7387 26581
rect 7283 26478 7387 26535
rect 7283 26432 7312 26478
rect 7358 26432 7387 26478
rect 7283 26375 7387 26432
rect 7283 26329 7312 26375
rect 7358 26329 7387 26375
rect 7283 26272 7387 26329
rect 7283 26226 7312 26272
rect 7358 26226 7387 26272
rect 7283 26169 7387 26226
rect 7283 26123 7312 26169
rect 7358 26123 7387 26169
rect 7283 26065 7387 26123
rect 7283 26019 7312 26065
rect 7358 26019 7387 26065
rect 7283 26006 7387 26019
rect 7527 26993 7631 27006
rect 7527 26947 7556 26993
rect 7602 26947 7631 26993
rect 7527 26890 7631 26947
rect 7527 26844 7556 26890
rect 7602 26844 7631 26890
rect 7527 26787 7631 26844
rect 7527 26741 7556 26787
rect 7602 26741 7631 26787
rect 7527 26684 7631 26741
rect 7527 26638 7556 26684
rect 7602 26638 7631 26684
rect 7527 26581 7631 26638
rect 7527 26535 7556 26581
rect 7602 26535 7631 26581
rect 7527 26478 7631 26535
rect 7527 26432 7556 26478
rect 7602 26432 7631 26478
rect 7527 26375 7631 26432
rect 7527 26329 7556 26375
rect 7602 26329 7631 26375
rect 7527 26272 7631 26329
rect 7527 26226 7556 26272
rect 7602 26226 7631 26272
rect 7527 26169 7631 26226
rect 7527 26123 7556 26169
rect 7602 26123 7631 26169
rect 7527 26065 7631 26123
rect 7527 26019 7556 26065
rect 7602 26019 7631 26065
rect 7527 26006 7631 26019
rect 7771 26993 7875 27006
rect 7771 26947 7800 26993
rect 7846 26947 7875 26993
rect 7771 26890 7875 26947
rect 7771 26844 7800 26890
rect 7846 26844 7875 26890
rect 7771 26787 7875 26844
rect 7771 26741 7800 26787
rect 7846 26741 7875 26787
rect 7771 26684 7875 26741
rect 7771 26638 7800 26684
rect 7846 26638 7875 26684
rect 7771 26581 7875 26638
rect 7771 26535 7800 26581
rect 7846 26535 7875 26581
rect 7771 26478 7875 26535
rect 7771 26432 7800 26478
rect 7846 26432 7875 26478
rect 7771 26375 7875 26432
rect 7771 26329 7800 26375
rect 7846 26329 7875 26375
rect 7771 26272 7875 26329
rect 7771 26226 7800 26272
rect 7846 26226 7875 26272
rect 7771 26169 7875 26226
rect 7771 26123 7800 26169
rect 7846 26123 7875 26169
rect 7771 26065 7875 26123
rect 7771 26019 7800 26065
rect 7846 26019 7875 26065
rect 7771 26006 7875 26019
rect 8015 26993 8103 27006
rect 8015 26947 8044 26993
rect 8090 26947 8103 26993
rect 8015 26890 8103 26947
rect 8015 26844 8044 26890
rect 8090 26844 8103 26890
rect 8015 26787 8103 26844
rect 8015 26741 8044 26787
rect 8090 26741 8103 26787
rect 8015 26684 8103 26741
rect 8015 26638 8044 26684
rect 8090 26638 8103 26684
rect 8015 26581 8103 26638
rect 8015 26535 8044 26581
rect 8090 26535 8103 26581
rect 8015 26478 8103 26535
rect 8015 26432 8044 26478
rect 8090 26432 8103 26478
rect 8015 26375 8103 26432
rect 8015 26329 8044 26375
rect 8090 26329 8103 26375
rect 8015 26272 8103 26329
rect 8015 26226 8044 26272
rect 8090 26226 8103 26272
rect 8015 26169 8103 26226
rect 8015 26123 8044 26169
rect 8090 26123 8103 26169
rect 8015 26065 8103 26123
rect 8015 26019 8044 26065
rect 8090 26019 8103 26065
rect 8015 26006 8103 26019
<< mvpdiff >>
rect 2577 28904 2665 28917
rect 2577 28858 2590 28904
rect 2636 28858 2665 28904
rect 2577 28801 2665 28858
rect 2577 28755 2590 28801
rect 2636 28755 2665 28801
rect 2577 28698 2665 28755
rect 2577 28652 2590 28698
rect 2636 28652 2665 28698
rect 2577 28595 2665 28652
rect 2577 28549 2590 28595
rect 2636 28549 2665 28595
rect 2577 28492 2665 28549
rect 2577 28446 2590 28492
rect 2636 28446 2665 28492
rect 2577 28389 2665 28446
rect 2577 28343 2590 28389
rect 2636 28343 2665 28389
rect 2577 28286 2665 28343
rect 2577 28240 2590 28286
rect 2636 28240 2665 28286
rect 2577 28183 2665 28240
rect 2577 28137 2590 28183
rect 2636 28137 2665 28183
rect 2577 28080 2665 28137
rect 2577 28034 2590 28080
rect 2636 28034 2665 28080
rect 2577 27976 2665 28034
rect 2577 27930 2590 27976
rect 2636 27930 2665 27976
rect 2577 27917 2665 27930
rect 2805 28904 2909 28917
rect 2805 28858 2834 28904
rect 2880 28858 2909 28904
rect 2805 28801 2909 28858
rect 2805 28755 2834 28801
rect 2880 28755 2909 28801
rect 2805 28698 2909 28755
rect 2805 28652 2834 28698
rect 2880 28652 2909 28698
rect 2805 28595 2909 28652
rect 2805 28549 2834 28595
rect 2880 28549 2909 28595
rect 2805 28492 2909 28549
rect 2805 28446 2834 28492
rect 2880 28446 2909 28492
rect 2805 28389 2909 28446
rect 2805 28343 2834 28389
rect 2880 28343 2909 28389
rect 2805 28286 2909 28343
rect 2805 28240 2834 28286
rect 2880 28240 2909 28286
rect 2805 28183 2909 28240
rect 2805 28137 2834 28183
rect 2880 28137 2909 28183
rect 2805 28080 2909 28137
rect 2805 28034 2834 28080
rect 2880 28034 2909 28080
rect 2805 27976 2909 28034
rect 2805 27930 2834 27976
rect 2880 27930 2909 27976
rect 2805 27917 2909 27930
rect 3049 28904 3153 28917
rect 3049 28858 3078 28904
rect 3124 28858 3153 28904
rect 3049 28801 3153 28858
rect 3049 28755 3078 28801
rect 3124 28755 3153 28801
rect 3049 28698 3153 28755
rect 3049 28652 3078 28698
rect 3124 28652 3153 28698
rect 3049 28595 3153 28652
rect 3049 28549 3078 28595
rect 3124 28549 3153 28595
rect 3049 28492 3153 28549
rect 3049 28446 3078 28492
rect 3124 28446 3153 28492
rect 3049 28389 3153 28446
rect 3049 28343 3078 28389
rect 3124 28343 3153 28389
rect 3049 28286 3153 28343
rect 3049 28240 3078 28286
rect 3124 28240 3153 28286
rect 3049 28183 3153 28240
rect 3049 28137 3078 28183
rect 3124 28137 3153 28183
rect 3049 28080 3153 28137
rect 3049 28034 3078 28080
rect 3124 28034 3153 28080
rect 3049 27976 3153 28034
rect 3049 27930 3078 27976
rect 3124 27930 3153 27976
rect 3049 27917 3153 27930
rect 3293 28904 3397 28917
rect 3293 28858 3322 28904
rect 3368 28858 3397 28904
rect 3293 28801 3397 28858
rect 3293 28755 3322 28801
rect 3368 28755 3397 28801
rect 3293 28698 3397 28755
rect 3293 28652 3322 28698
rect 3368 28652 3397 28698
rect 3293 28595 3397 28652
rect 3293 28549 3322 28595
rect 3368 28549 3397 28595
rect 3293 28492 3397 28549
rect 3293 28446 3322 28492
rect 3368 28446 3397 28492
rect 3293 28389 3397 28446
rect 3293 28343 3322 28389
rect 3368 28343 3397 28389
rect 3293 28286 3397 28343
rect 3293 28240 3322 28286
rect 3368 28240 3397 28286
rect 3293 28183 3397 28240
rect 3293 28137 3322 28183
rect 3368 28137 3397 28183
rect 3293 28080 3397 28137
rect 3293 28034 3322 28080
rect 3368 28034 3397 28080
rect 3293 27976 3397 28034
rect 3293 27930 3322 27976
rect 3368 27930 3397 27976
rect 3293 27917 3397 27930
rect 3537 28904 3641 28917
rect 3537 28858 3566 28904
rect 3612 28858 3641 28904
rect 3537 28801 3641 28858
rect 3537 28755 3566 28801
rect 3612 28755 3641 28801
rect 3537 28698 3641 28755
rect 3537 28652 3566 28698
rect 3612 28652 3641 28698
rect 3537 28595 3641 28652
rect 3537 28549 3566 28595
rect 3612 28549 3641 28595
rect 3537 28492 3641 28549
rect 3537 28446 3566 28492
rect 3612 28446 3641 28492
rect 3537 28389 3641 28446
rect 3537 28343 3566 28389
rect 3612 28343 3641 28389
rect 3537 28286 3641 28343
rect 3537 28240 3566 28286
rect 3612 28240 3641 28286
rect 3537 28183 3641 28240
rect 3537 28137 3566 28183
rect 3612 28137 3641 28183
rect 3537 28080 3641 28137
rect 3537 28034 3566 28080
rect 3612 28034 3641 28080
rect 3537 27976 3641 28034
rect 3537 27930 3566 27976
rect 3612 27930 3641 27976
rect 3537 27917 3641 27930
rect 3781 28904 3885 28917
rect 3781 28858 3810 28904
rect 3856 28858 3885 28904
rect 3781 28801 3885 28858
rect 3781 28755 3810 28801
rect 3856 28755 3885 28801
rect 3781 28698 3885 28755
rect 3781 28652 3810 28698
rect 3856 28652 3885 28698
rect 3781 28595 3885 28652
rect 3781 28549 3810 28595
rect 3856 28549 3885 28595
rect 3781 28492 3885 28549
rect 3781 28446 3810 28492
rect 3856 28446 3885 28492
rect 3781 28389 3885 28446
rect 3781 28343 3810 28389
rect 3856 28343 3885 28389
rect 3781 28286 3885 28343
rect 3781 28240 3810 28286
rect 3856 28240 3885 28286
rect 3781 28183 3885 28240
rect 3781 28137 3810 28183
rect 3856 28137 3885 28183
rect 3781 28080 3885 28137
rect 3781 28034 3810 28080
rect 3856 28034 3885 28080
rect 3781 27976 3885 28034
rect 3781 27930 3810 27976
rect 3856 27930 3885 27976
rect 3781 27917 3885 27930
rect 4025 28904 4129 28917
rect 4025 28858 4054 28904
rect 4100 28858 4129 28904
rect 4025 28801 4129 28858
rect 4025 28755 4054 28801
rect 4100 28755 4129 28801
rect 4025 28698 4129 28755
rect 4025 28652 4054 28698
rect 4100 28652 4129 28698
rect 4025 28595 4129 28652
rect 4025 28549 4054 28595
rect 4100 28549 4129 28595
rect 4025 28492 4129 28549
rect 4025 28446 4054 28492
rect 4100 28446 4129 28492
rect 4025 28389 4129 28446
rect 4025 28343 4054 28389
rect 4100 28343 4129 28389
rect 4025 28286 4129 28343
rect 4025 28240 4054 28286
rect 4100 28240 4129 28286
rect 4025 28183 4129 28240
rect 4025 28137 4054 28183
rect 4100 28137 4129 28183
rect 4025 28080 4129 28137
rect 4025 28034 4054 28080
rect 4100 28034 4129 28080
rect 4025 27976 4129 28034
rect 4025 27930 4054 27976
rect 4100 27930 4129 27976
rect 4025 27917 4129 27930
rect 4269 28904 4357 28917
rect 4269 28858 4298 28904
rect 4344 28858 4357 28904
rect 4269 28801 4357 28858
rect 4269 28755 4298 28801
rect 4344 28755 4357 28801
rect 4269 28698 4357 28755
rect 4269 28652 4298 28698
rect 4344 28652 4357 28698
rect 4269 28595 4357 28652
rect 4269 28549 4298 28595
rect 4344 28549 4357 28595
rect 4269 28492 4357 28549
rect 4269 28446 4298 28492
rect 4344 28446 4357 28492
rect 4269 28389 4357 28446
rect 4269 28343 4298 28389
rect 4344 28343 4357 28389
rect 4269 28286 4357 28343
rect 4269 28240 4298 28286
rect 4344 28240 4357 28286
rect 4269 28183 4357 28240
rect 4269 28137 4298 28183
rect 4344 28137 4357 28183
rect 4269 28080 4357 28137
rect 4269 28034 4298 28080
rect 4344 28034 4357 28080
rect 4269 27976 4357 28034
rect 4269 27930 4298 27976
rect 4344 27930 4357 27976
rect 4269 27917 4357 27930
rect 4457 28904 4545 28917
rect 4457 28858 4470 28904
rect 4516 28858 4545 28904
rect 4457 28801 4545 28858
rect 4457 28755 4470 28801
rect 4516 28755 4545 28801
rect 4457 28698 4545 28755
rect 4457 28652 4470 28698
rect 4516 28652 4545 28698
rect 4457 28595 4545 28652
rect 4457 28549 4470 28595
rect 4516 28549 4545 28595
rect 4457 28492 4545 28549
rect 4457 28446 4470 28492
rect 4516 28446 4545 28492
rect 4457 28389 4545 28446
rect 4457 28343 4470 28389
rect 4516 28343 4545 28389
rect 4457 28286 4545 28343
rect 4457 28240 4470 28286
rect 4516 28240 4545 28286
rect 4457 28183 4545 28240
rect 4457 28137 4470 28183
rect 4516 28137 4545 28183
rect 4457 28080 4545 28137
rect 4457 28034 4470 28080
rect 4516 28034 4545 28080
rect 4457 27976 4545 28034
rect 4457 27930 4470 27976
rect 4516 27930 4545 27976
rect 4457 27917 4545 27930
rect 4685 28904 4789 28917
rect 4685 28858 4714 28904
rect 4760 28858 4789 28904
rect 4685 28801 4789 28858
rect 4685 28755 4714 28801
rect 4760 28755 4789 28801
rect 4685 28698 4789 28755
rect 4685 28652 4714 28698
rect 4760 28652 4789 28698
rect 4685 28595 4789 28652
rect 4685 28549 4714 28595
rect 4760 28549 4789 28595
rect 4685 28492 4789 28549
rect 4685 28446 4714 28492
rect 4760 28446 4789 28492
rect 4685 28389 4789 28446
rect 4685 28343 4714 28389
rect 4760 28343 4789 28389
rect 4685 28286 4789 28343
rect 4685 28240 4714 28286
rect 4760 28240 4789 28286
rect 4685 28183 4789 28240
rect 4685 28137 4714 28183
rect 4760 28137 4789 28183
rect 4685 28080 4789 28137
rect 4685 28034 4714 28080
rect 4760 28034 4789 28080
rect 4685 27976 4789 28034
rect 4685 27930 4714 27976
rect 4760 27930 4789 27976
rect 4685 27917 4789 27930
rect 4929 28904 5033 28917
rect 4929 28858 4958 28904
rect 5004 28858 5033 28904
rect 4929 28801 5033 28858
rect 4929 28755 4958 28801
rect 5004 28755 5033 28801
rect 4929 28698 5033 28755
rect 4929 28652 4958 28698
rect 5004 28652 5033 28698
rect 4929 28595 5033 28652
rect 4929 28549 4958 28595
rect 5004 28549 5033 28595
rect 4929 28492 5033 28549
rect 4929 28446 4958 28492
rect 5004 28446 5033 28492
rect 4929 28389 5033 28446
rect 4929 28343 4958 28389
rect 5004 28343 5033 28389
rect 4929 28286 5033 28343
rect 4929 28240 4958 28286
rect 5004 28240 5033 28286
rect 4929 28183 5033 28240
rect 4929 28137 4958 28183
rect 5004 28137 5033 28183
rect 4929 28080 5033 28137
rect 4929 28034 4958 28080
rect 5004 28034 5033 28080
rect 4929 27976 5033 28034
rect 4929 27930 4958 27976
rect 5004 27930 5033 27976
rect 4929 27917 5033 27930
rect 5173 28904 5277 28917
rect 5173 28858 5202 28904
rect 5248 28858 5277 28904
rect 5173 28801 5277 28858
rect 5173 28755 5202 28801
rect 5248 28755 5277 28801
rect 5173 28698 5277 28755
rect 5173 28652 5202 28698
rect 5248 28652 5277 28698
rect 5173 28595 5277 28652
rect 5173 28549 5202 28595
rect 5248 28549 5277 28595
rect 5173 28492 5277 28549
rect 5173 28446 5202 28492
rect 5248 28446 5277 28492
rect 5173 28389 5277 28446
rect 5173 28343 5202 28389
rect 5248 28343 5277 28389
rect 5173 28286 5277 28343
rect 5173 28240 5202 28286
rect 5248 28240 5277 28286
rect 5173 28183 5277 28240
rect 5173 28137 5202 28183
rect 5248 28137 5277 28183
rect 5173 28080 5277 28137
rect 5173 28034 5202 28080
rect 5248 28034 5277 28080
rect 5173 27976 5277 28034
rect 5173 27930 5202 27976
rect 5248 27930 5277 27976
rect 5173 27917 5277 27930
rect 5417 28904 5521 28917
rect 5417 28858 5446 28904
rect 5492 28858 5521 28904
rect 5417 28801 5521 28858
rect 5417 28755 5446 28801
rect 5492 28755 5521 28801
rect 5417 28698 5521 28755
rect 5417 28652 5446 28698
rect 5492 28652 5521 28698
rect 5417 28595 5521 28652
rect 5417 28549 5446 28595
rect 5492 28549 5521 28595
rect 5417 28492 5521 28549
rect 5417 28446 5446 28492
rect 5492 28446 5521 28492
rect 5417 28389 5521 28446
rect 5417 28343 5446 28389
rect 5492 28343 5521 28389
rect 5417 28286 5521 28343
rect 5417 28240 5446 28286
rect 5492 28240 5521 28286
rect 5417 28183 5521 28240
rect 5417 28137 5446 28183
rect 5492 28137 5521 28183
rect 5417 28080 5521 28137
rect 5417 28034 5446 28080
rect 5492 28034 5521 28080
rect 5417 27976 5521 28034
rect 5417 27930 5446 27976
rect 5492 27930 5521 27976
rect 5417 27917 5521 27930
rect 5661 28904 5765 28917
rect 5661 28858 5690 28904
rect 5736 28858 5765 28904
rect 5661 28801 5765 28858
rect 5661 28755 5690 28801
rect 5736 28755 5765 28801
rect 5661 28698 5765 28755
rect 5661 28652 5690 28698
rect 5736 28652 5765 28698
rect 5661 28595 5765 28652
rect 5661 28549 5690 28595
rect 5736 28549 5765 28595
rect 5661 28492 5765 28549
rect 5661 28446 5690 28492
rect 5736 28446 5765 28492
rect 5661 28389 5765 28446
rect 5661 28343 5690 28389
rect 5736 28343 5765 28389
rect 5661 28286 5765 28343
rect 5661 28240 5690 28286
rect 5736 28240 5765 28286
rect 5661 28183 5765 28240
rect 5661 28137 5690 28183
rect 5736 28137 5765 28183
rect 5661 28080 5765 28137
rect 5661 28034 5690 28080
rect 5736 28034 5765 28080
rect 5661 27976 5765 28034
rect 5661 27930 5690 27976
rect 5736 27930 5765 27976
rect 5661 27917 5765 27930
rect 5905 28904 6009 28917
rect 5905 28858 5934 28904
rect 5980 28858 6009 28904
rect 5905 28801 6009 28858
rect 5905 28755 5934 28801
rect 5980 28755 6009 28801
rect 5905 28698 6009 28755
rect 5905 28652 5934 28698
rect 5980 28652 6009 28698
rect 5905 28595 6009 28652
rect 5905 28549 5934 28595
rect 5980 28549 6009 28595
rect 5905 28492 6009 28549
rect 5905 28446 5934 28492
rect 5980 28446 6009 28492
rect 5905 28389 6009 28446
rect 5905 28343 5934 28389
rect 5980 28343 6009 28389
rect 5905 28286 6009 28343
rect 5905 28240 5934 28286
rect 5980 28240 6009 28286
rect 5905 28183 6009 28240
rect 5905 28137 5934 28183
rect 5980 28137 6009 28183
rect 5905 28080 6009 28137
rect 5905 28034 5934 28080
rect 5980 28034 6009 28080
rect 5905 27976 6009 28034
rect 5905 27930 5934 27976
rect 5980 27930 6009 27976
rect 5905 27917 6009 27930
rect 6149 28904 6253 28917
rect 6149 28858 6178 28904
rect 6224 28858 6253 28904
rect 6149 28801 6253 28858
rect 6149 28755 6178 28801
rect 6224 28755 6253 28801
rect 6149 28698 6253 28755
rect 6149 28652 6178 28698
rect 6224 28652 6253 28698
rect 6149 28595 6253 28652
rect 6149 28549 6178 28595
rect 6224 28549 6253 28595
rect 6149 28492 6253 28549
rect 6149 28446 6178 28492
rect 6224 28446 6253 28492
rect 6149 28389 6253 28446
rect 6149 28343 6178 28389
rect 6224 28343 6253 28389
rect 6149 28286 6253 28343
rect 6149 28240 6178 28286
rect 6224 28240 6253 28286
rect 6149 28183 6253 28240
rect 6149 28137 6178 28183
rect 6224 28137 6253 28183
rect 6149 28080 6253 28137
rect 6149 28034 6178 28080
rect 6224 28034 6253 28080
rect 6149 27976 6253 28034
rect 6149 27930 6178 27976
rect 6224 27930 6253 27976
rect 6149 27917 6253 27930
rect 6393 28904 6497 28917
rect 6393 28858 6422 28904
rect 6468 28858 6497 28904
rect 6393 28801 6497 28858
rect 6393 28755 6422 28801
rect 6468 28755 6497 28801
rect 6393 28698 6497 28755
rect 6393 28652 6422 28698
rect 6468 28652 6497 28698
rect 6393 28595 6497 28652
rect 6393 28549 6422 28595
rect 6468 28549 6497 28595
rect 6393 28492 6497 28549
rect 6393 28446 6422 28492
rect 6468 28446 6497 28492
rect 6393 28389 6497 28446
rect 6393 28343 6422 28389
rect 6468 28343 6497 28389
rect 6393 28286 6497 28343
rect 6393 28240 6422 28286
rect 6468 28240 6497 28286
rect 6393 28183 6497 28240
rect 6393 28137 6422 28183
rect 6468 28137 6497 28183
rect 6393 28080 6497 28137
rect 6393 28034 6422 28080
rect 6468 28034 6497 28080
rect 6393 27976 6497 28034
rect 6393 27930 6422 27976
rect 6468 27930 6497 27976
rect 6393 27917 6497 27930
rect 6637 28904 6741 28917
rect 6637 28858 6666 28904
rect 6712 28858 6741 28904
rect 6637 28801 6741 28858
rect 6637 28755 6666 28801
rect 6712 28755 6741 28801
rect 6637 28698 6741 28755
rect 6637 28652 6666 28698
rect 6712 28652 6741 28698
rect 6637 28595 6741 28652
rect 6637 28549 6666 28595
rect 6712 28549 6741 28595
rect 6637 28492 6741 28549
rect 6637 28446 6666 28492
rect 6712 28446 6741 28492
rect 6637 28389 6741 28446
rect 6637 28343 6666 28389
rect 6712 28343 6741 28389
rect 6637 28286 6741 28343
rect 6637 28240 6666 28286
rect 6712 28240 6741 28286
rect 6637 28183 6741 28240
rect 6637 28137 6666 28183
rect 6712 28137 6741 28183
rect 6637 28080 6741 28137
rect 6637 28034 6666 28080
rect 6712 28034 6741 28080
rect 6637 27976 6741 28034
rect 6637 27930 6666 27976
rect 6712 27930 6741 27976
rect 6637 27917 6741 27930
rect 6881 28904 6985 28917
rect 6881 28858 6910 28904
rect 6956 28858 6985 28904
rect 6881 28801 6985 28858
rect 6881 28755 6910 28801
rect 6956 28755 6985 28801
rect 6881 28698 6985 28755
rect 6881 28652 6910 28698
rect 6956 28652 6985 28698
rect 6881 28595 6985 28652
rect 6881 28549 6910 28595
rect 6956 28549 6985 28595
rect 6881 28492 6985 28549
rect 6881 28446 6910 28492
rect 6956 28446 6985 28492
rect 6881 28389 6985 28446
rect 6881 28343 6910 28389
rect 6956 28343 6985 28389
rect 6881 28286 6985 28343
rect 6881 28240 6910 28286
rect 6956 28240 6985 28286
rect 6881 28183 6985 28240
rect 6881 28137 6910 28183
rect 6956 28137 6985 28183
rect 6881 28080 6985 28137
rect 6881 28034 6910 28080
rect 6956 28034 6985 28080
rect 6881 27976 6985 28034
rect 6881 27930 6910 27976
rect 6956 27930 6985 27976
rect 6881 27917 6985 27930
rect 7125 28904 7229 28917
rect 7125 28858 7154 28904
rect 7200 28858 7229 28904
rect 7125 28801 7229 28858
rect 7125 28755 7154 28801
rect 7200 28755 7229 28801
rect 7125 28698 7229 28755
rect 7125 28652 7154 28698
rect 7200 28652 7229 28698
rect 7125 28595 7229 28652
rect 7125 28549 7154 28595
rect 7200 28549 7229 28595
rect 7125 28492 7229 28549
rect 7125 28446 7154 28492
rect 7200 28446 7229 28492
rect 7125 28389 7229 28446
rect 7125 28343 7154 28389
rect 7200 28343 7229 28389
rect 7125 28286 7229 28343
rect 7125 28240 7154 28286
rect 7200 28240 7229 28286
rect 7125 28183 7229 28240
rect 7125 28137 7154 28183
rect 7200 28137 7229 28183
rect 7125 28080 7229 28137
rect 7125 28034 7154 28080
rect 7200 28034 7229 28080
rect 7125 27976 7229 28034
rect 7125 27930 7154 27976
rect 7200 27930 7229 27976
rect 7125 27917 7229 27930
rect 7369 28904 7473 28917
rect 7369 28858 7398 28904
rect 7444 28858 7473 28904
rect 7369 28801 7473 28858
rect 7369 28755 7398 28801
rect 7444 28755 7473 28801
rect 7369 28698 7473 28755
rect 7369 28652 7398 28698
rect 7444 28652 7473 28698
rect 7369 28595 7473 28652
rect 7369 28549 7398 28595
rect 7444 28549 7473 28595
rect 7369 28492 7473 28549
rect 7369 28446 7398 28492
rect 7444 28446 7473 28492
rect 7369 28389 7473 28446
rect 7369 28343 7398 28389
rect 7444 28343 7473 28389
rect 7369 28286 7473 28343
rect 7369 28240 7398 28286
rect 7444 28240 7473 28286
rect 7369 28183 7473 28240
rect 7369 28137 7398 28183
rect 7444 28137 7473 28183
rect 7369 28080 7473 28137
rect 7369 28034 7398 28080
rect 7444 28034 7473 28080
rect 7369 27976 7473 28034
rect 7369 27930 7398 27976
rect 7444 27930 7473 27976
rect 7369 27917 7473 27930
rect 7613 28904 7717 28917
rect 7613 28858 7642 28904
rect 7688 28858 7717 28904
rect 7613 28801 7717 28858
rect 7613 28755 7642 28801
rect 7688 28755 7717 28801
rect 7613 28698 7717 28755
rect 7613 28652 7642 28698
rect 7688 28652 7717 28698
rect 7613 28595 7717 28652
rect 7613 28549 7642 28595
rect 7688 28549 7717 28595
rect 7613 28492 7717 28549
rect 7613 28446 7642 28492
rect 7688 28446 7717 28492
rect 7613 28389 7717 28446
rect 7613 28343 7642 28389
rect 7688 28343 7717 28389
rect 7613 28286 7717 28343
rect 7613 28240 7642 28286
rect 7688 28240 7717 28286
rect 7613 28183 7717 28240
rect 7613 28137 7642 28183
rect 7688 28137 7717 28183
rect 7613 28080 7717 28137
rect 7613 28034 7642 28080
rect 7688 28034 7717 28080
rect 7613 27976 7717 28034
rect 7613 27930 7642 27976
rect 7688 27930 7717 27976
rect 7613 27917 7717 27930
rect 7857 28904 7961 28917
rect 7857 28858 7886 28904
rect 7932 28858 7961 28904
rect 7857 28801 7961 28858
rect 7857 28755 7886 28801
rect 7932 28755 7961 28801
rect 7857 28698 7961 28755
rect 7857 28652 7886 28698
rect 7932 28652 7961 28698
rect 7857 28595 7961 28652
rect 7857 28549 7886 28595
rect 7932 28549 7961 28595
rect 7857 28492 7961 28549
rect 7857 28446 7886 28492
rect 7932 28446 7961 28492
rect 7857 28389 7961 28446
rect 7857 28343 7886 28389
rect 7932 28343 7961 28389
rect 7857 28286 7961 28343
rect 7857 28240 7886 28286
rect 7932 28240 7961 28286
rect 7857 28183 7961 28240
rect 7857 28137 7886 28183
rect 7932 28137 7961 28183
rect 7857 28080 7961 28137
rect 7857 28034 7886 28080
rect 7932 28034 7961 28080
rect 7857 27976 7961 28034
rect 7857 27930 7886 27976
rect 7932 27930 7961 27976
rect 7857 27917 7961 27930
rect 8101 28904 8205 28917
rect 8101 28858 8130 28904
rect 8176 28858 8205 28904
rect 8101 28801 8205 28858
rect 8101 28755 8130 28801
rect 8176 28755 8205 28801
rect 8101 28698 8205 28755
rect 8101 28652 8130 28698
rect 8176 28652 8205 28698
rect 8101 28595 8205 28652
rect 8101 28549 8130 28595
rect 8176 28549 8205 28595
rect 8101 28492 8205 28549
rect 8101 28446 8130 28492
rect 8176 28446 8205 28492
rect 8101 28389 8205 28446
rect 8101 28343 8130 28389
rect 8176 28343 8205 28389
rect 8101 28286 8205 28343
rect 8101 28240 8130 28286
rect 8176 28240 8205 28286
rect 8101 28183 8205 28240
rect 8101 28137 8130 28183
rect 8176 28137 8205 28183
rect 8101 28080 8205 28137
rect 8101 28034 8130 28080
rect 8176 28034 8205 28080
rect 8101 27976 8205 28034
rect 8101 27930 8130 27976
rect 8176 27930 8205 27976
rect 8101 27917 8205 27930
rect 8345 28904 8449 28917
rect 8345 28858 8374 28904
rect 8420 28858 8449 28904
rect 8345 28801 8449 28858
rect 8345 28755 8374 28801
rect 8420 28755 8449 28801
rect 8345 28698 8449 28755
rect 8345 28652 8374 28698
rect 8420 28652 8449 28698
rect 8345 28595 8449 28652
rect 8345 28549 8374 28595
rect 8420 28549 8449 28595
rect 8345 28492 8449 28549
rect 8345 28446 8374 28492
rect 8420 28446 8449 28492
rect 8345 28389 8449 28446
rect 8345 28343 8374 28389
rect 8420 28343 8449 28389
rect 8345 28286 8449 28343
rect 8345 28240 8374 28286
rect 8420 28240 8449 28286
rect 8345 28183 8449 28240
rect 8345 28137 8374 28183
rect 8420 28137 8449 28183
rect 8345 28080 8449 28137
rect 8345 28034 8374 28080
rect 8420 28034 8449 28080
rect 8345 27976 8449 28034
rect 8345 27930 8374 27976
rect 8420 27930 8449 27976
rect 8345 27917 8449 27930
rect 8589 28904 8693 28917
rect 8589 28858 8618 28904
rect 8664 28858 8693 28904
rect 8589 28801 8693 28858
rect 8589 28755 8618 28801
rect 8664 28755 8693 28801
rect 8589 28698 8693 28755
rect 8589 28652 8618 28698
rect 8664 28652 8693 28698
rect 8589 28595 8693 28652
rect 8589 28549 8618 28595
rect 8664 28549 8693 28595
rect 8589 28492 8693 28549
rect 8589 28446 8618 28492
rect 8664 28446 8693 28492
rect 8589 28389 8693 28446
rect 8589 28343 8618 28389
rect 8664 28343 8693 28389
rect 8589 28286 8693 28343
rect 8589 28240 8618 28286
rect 8664 28240 8693 28286
rect 8589 28183 8693 28240
rect 8589 28137 8618 28183
rect 8664 28137 8693 28183
rect 8589 28080 8693 28137
rect 8589 28034 8618 28080
rect 8664 28034 8693 28080
rect 8589 27976 8693 28034
rect 8589 27930 8618 27976
rect 8664 27930 8693 27976
rect 8589 27917 8693 27930
rect 8833 28904 8937 28917
rect 8833 28858 8862 28904
rect 8908 28858 8937 28904
rect 8833 28801 8937 28858
rect 8833 28755 8862 28801
rect 8908 28755 8937 28801
rect 8833 28698 8937 28755
rect 8833 28652 8862 28698
rect 8908 28652 8937 28698
rect 8833 28595 8937 28652
rect 8833 28549 8862 28595
rect 8908 28549 8937 28595
rect 8833 28492 8937 28549
rect 8833 28446 8862 28492
rect 8908 28446 8937 28492
rect 8833 28389 8937 28446
rect 8833 28343 8862 28389
rect 8908 28343 8937 28389
rect 8833 28286 8937 28343
rect 8833 28240 8862 28286
rect 8908 28240 8937 28286
rect 8833 28183 8937 28240
rect 8833 28137 8862 28183
rect 8908 28137 8937 28183
rect 8833 28080 8937 28137
rect 8833 28034 8862 28080
rect 8908 28034 8937 28080
rect 8833 27976 8937 28034
rect 8833 27930 8862 27976
rect 8908 27930 8937 27976
rect 8833 27917 8937 27930
rect 9077 28904 9181 28917
rect 9077 28858 9106 28904
rect 9152 28858 9181 28904
rect 9077 28801 9181 28858
rect 9077 28755 9106 28801
rect 9152 28755 9181 28801
rect 9077 28698 9181 28755
rect 9077 28652 9106 28698
rect 9152 28652 9181 28698
rect 9077 28595 9181 28652
rect 9077 28549 9106 28595
rect 9152 28549 9181 28595
rect 9077 28492 9181 28549
rect 9077 28446 9106 28492
rect 9152 28446 9181 28492
rect 9077 28389 9181 28446
rect 9077 28343 9106 28389
rect 9152 28343 9181 28389
rect 9077 28286 9181 28343
rect 9077 28240 9106 28286
rect 9152 28240 9181 28286
rect 9077 28183 9181 28240
rect 9077 28137 9106 28183
rect 9152 28137 9181 28183
rect 9077 28080 9181 28137
rect 9077 28034 9106 28080
rect 9152 28034 9181 28080
rect 9077 27976 9181 28034
rect 9077 27930 9106 27976
rect 9152 27930 9181 27976
rect 9077 27917 9181 27930
rect 9321 28904 9425 28917
rect 9321 28858 9350 28904
rect 9396 28858 9425 28904
rect 9321 28801 9425 28858
rect 9321 28755 9350 28801
rect 9396 28755 9425 28801
rect 9321 28698 9425 28755
rect 9321 28652 9350 28698
rect 9396 28652 9425 28698
rect 9321 28595 9425 28652
rect 9321 28549 9350 28595
rect 9396 28549 9425 28595
rect 9321 28492 9425 28549
rect 9321 28446 9350 28492
rect 9396 28446 9425 28492
rect 9321 28389 9425 28446
rect 9321 28343 9350 28389
rect 9396 28343 9425 28389
rect 9321 28286 9425 28343
rect 9321 28240 9350 28286
rect 9396 28240 9425 28286
rect 9321 28183 9425 28240
rect 9321 28137 9350 28183
rect 9396 28137 9425 28183
rect 9321 28080 9425 28137
rect 9321 28034 9350 28080
rect 9396 28034 9425 28080
rect 9321 27976 9425 28034
rect 9321 27930 9350 27976
rect 9396 27930 9425 27976
rect 9321 27917 9425 27930
rect 9565 28904 9669 28917
rect 9565 28858 9594 28904
rect 9640 28858 9669 28904
rect 9565 28801 9669 28858
rect 9565 28755 9594 28801
rect 9640 28755 9669 28801
rect 9565 28698 9669 28755
rect 9565 28652 9594 28698
rect 9640 28652 9669 28698
rect 9565 28595 9669 28652
rect 9565 28549 9594 28595
rect 9640 28549 9669 28595
rect 9565 28492 9669 28549
rect 9565 28446 9594 28492
rect 9640 28446 9669 28492
rect 9565 28389 9669 28446
rect 9565 28343 9594 28389
rect 9640 28343 9669 28389
rect 9565 28286 9669 28343
rect 9565 28240 9594 28286
rect 9640 28240 9669 28286
rect 9565 28183 9669 28240
rect 9565 28137 9594 28183
rect 9640 28137 9669 28183
rect 9565 28080 9669 28137
rect 9565 28034 9594 28080
rect 9640 28034 9669 28080
rect 9565 27976 9669 28034
rect 9565 27930 9594 27976
rect 9640 27930 9669 27976
rect 9565 27917 9669 27930
rect 9809 28904 9913 28917
rect 9809 28858 9838 28904
rect 9884 28858 9913 28904
rect 9809 28801 9913 28858
rect 9809 28755 9838 28801
rect 9884 28755 9913 28801
rect 9809 28698 9913 28755
rect 9809 28652 9838 28698
rect 9884 28652 9913 28698
rect 9809 28595 9913 28652
rect 9809 28549 9838 28595
rect 9884 28549 9913 28595
rect 9809 28492 9913 28549
rect 9809 28446 9838 28492
rect 9884 28446 9913 28492
rect 9809 28389 9913 28446
rect 9809 28343 9838 28389
rect 9884 28343 9913 28389
rect 9809 28286 9913 28343
rect 9809 28240 9838 28286
rect 9884 28240 9913 28286
rect 9809 28183 9913 28240
rect 9809 28137 9838 28183
rect 9884 28137 9913 28183
rect 9809 28080 9913 28137
rect 9809 28034 9838 28080
rect 9884 28034 9913 28080
rect 9809 27976 9913 28034
rect 9809 27930 9838 27976
rect 9884 27930 9913 27976
rect 9809 27917 9913 27930
rect 10053 28904 10157 28917
rect 10053 28858 10082 28904
rect 10128 28858 10157 28904
rect 10053 28801 10157 28858
rect 10053 28755 10082 28801
rect 10128 28755 10157 28801
rect 10053 28698 10157 28755
rect 10053 28652 10082 28698
rect 10128 28652 10157 28698
rect 10053 28595 10157 28652
rect 10053 28549 10082 28595
rect 10128 28549 10157 28595
rect 10053 28492 10157 28549
rect 10053 28446 10082 28492
rect 10128 28446 10157 28492
rect 10053 28389 10157 28446
rect 10053 28343 10082 28389
rect 10128 28343 10157 28389
rect 10053 28286 10157 28343
rect 10053 28240 10082 28286
rect 10128 28240 10157 28286
rect 10053 28183 10157 28240
rect 10053 28137 10082 28183
rect 10128 28137 10157 28183
rect 10053 28080 10157 28137
rect 10053 28034 10082 28080
rect 10128 28034 10157 28080
rect 10053 27976 10157 28034
rect 10053 27930 10082 27976
rect 10128 27930 10157 27976
rect 10053 27917 10157 27930
rect 10297 28904 10385 28917
rect 10297 28858 10326 28904
rect 10372 28858 10385 28904
rect 10297 28801 10385 28858
rect 10297 28755 10326 28801
rect 10372 28755 10385 28801
rect 10297 28698 10385 28755
rect 10297 28652 10326 28698
rect 10372 28652 10385 28698
rect 10297 28595 10385 28652
rect 10297 28549 10326 28595
rect 10372 28549 10385 28595
rect 10297 28492 10385 28549
rect 10297 28446 10326 28492
rect 10372 28446 10385 28492
rect 10297 28389 10385 28446
rect 10297 28343 10326 28389
rect 10372 28343 10385 28389
rect 10297 28286 10385 28343
rect 10297 28240 10326 28286
rect 10372 28240 10385 28286
rect 10297 28183 10385 28240
rect 10297 28137 10326 28183
rect 10372 28137 10385 28183
rect 10297 28080 10385 28137
rect 10297 28034 10326 28080
rect 10372 28034 10385 28080
rect 10297 27976 10385 28034
rect 10297 27930 10326 27976
rect 10372 27930 10385 27976
rect 10297 27917 10385 27930
<< mvndiffc >>
rect 4054 26947 4100 26993
rect 4054 26844 4100 26890
rect 4054 26741 4100 26787
rect 4054 26638 4100 26684
rect 4054 26535 4100 26581
rect 4054 26432 4100 26478
rect 4054 26329 4100 26375
rect 4054 26226 4100 26272
rect 4054 26123 4100 26169
rect 4054 26019 4100 26065
rect 4298 26947 4344 26993
rect 4298 26844 4344 26890
rect 4298 26741 4344 26787
rect 4298 26638 4344 26684
rect 4298 26535 4344 26581
rect 4298 26432 4344 26478
rect 4298 26329 4344 26375
rect 4298 26226 4344 26272
rect 4298 26123 4344 26169
rect 4298 26019 4344 26065
rect 5116 26947 5162 26993
rect 5116 26844 5162 26890
rect 5116 26741 5162 26787
rect 5116 26638 5162 26684
rect 5116 26535 5162 26581
rect 5116 26432 5162 26478
rect 5116 26329 5162 26375
rect 5116 26226 5162 26272
rect 5116 26123 5162 26169
rect 5116 26019 5162 26065
rect 5360 26947 5406 26993
rect 5360 26844 5406 26890
rect 5360 26741 5406 26787
rect 5360 26638 5406 26684
rect 5360 26535 5406 26581
rect 5360 26432 5406 26478
rect 5360 26329 5406 26375
rect 5360 26226 5406 26272
rect 5360 26123 5406 26169
rect 5360 26019 5406 26065
rect 5604 26947 5650 26993
rect 5604 26844 5650 26890
rect 5604 26741 5650 26787
rect 5604 26638 5650 26684
rect 5604 26535 5650 26581
rect 5604 26432 5650 26478
rect 5604 26329 5650 26375
rect 5604 26226 5650 26272
rect 5604 26123 5650 26169
rect 5604 26019 5650 26065
rect 5848 26947 5894 26993
rect 5848 26844 5894 26890
rect 5848 26741 5894 26787
rect 5848 26638 5894 26684
rect 5848 26535 5894 26581
rect 5848 26432 5894 26478
rect 5848 26329 5894 26375
rect 5848 26226 5894 26272
rect 5848 26123 5894 26169
rect 5848 26019 5894 26065
rect 6092 26947 6138 26993
rect 6092 26844 6138 26890
rect 6092 26741 6138 26787
rect 6092 26638 6138 26684
rect 6092 26535 6138 26581
rect 6092 26432 6138 26478
rect 6092 26329 6138 26375
rect 6092 26226 6138 26272
rect 6092 26123 6138 26169
rect 6092 26019 6138 26065
rect 6336 26947 6382 26993
rect 6336 26844 6382 26890
rect 6336 26741 6382 26787
rect 6336 26638 6382 26684
rect 6336 26535 6382 26581
rect 6336 26432 6382 26478
rect 6336 26329 6382 26375
rect 6336 26226 6382 26272
rect 6336 26123 6382 26169
rect 6336 26019 6382 26065
rect 6580 26947 6626 26993
rect 6580 26844 6626 26890
rect 6580 26741 6626 26787
rect 6580 26638 6626 26684
rect 6580 26535 6626 26581
rect 6580 26432 6626 26478
rect 6580 26329 6626 26375
rect 6580 26226 6626 26272
rect 6580 26123 6626 26169
rect 6580 26019 6626 26065
rect 6824 26947 6870 26993
rect 6824 26844 6870 26890
rect 6824 26741 6870 26787
rect 6824 26638 6870 26684
rect 6824 26535 6870 26581
rect 6824 26432 6870 26478
rect 6824 26329 6870 26375
rect 6824 26226 6870 26272
rect 6824 26123 6870 26169
rect 6824 26019 6870 26065
rect 7068 26947 7114 26993
rect 7068 26844 7114 26890
rect 7068 26741 7114 26787
rect 7068 26638 7114 26684
rect 7068 26535 7114 26581
rect 7068 26432 7114 26478
rect 7068 26329 7114 26375
rect 7068 26226 7114 26272
rect 7068 26123 7114 26169
rect 7068 26019 7114 26065
rect 7312 26947 7358 26993
rect 7312 26844 7358 26890
rect 7312 26741 7358 26787
rect 7312 26638 7358 26684
rect 7312 26535 7358 26581
rect 7312 26432 7358 26478
rect 7312 26329 7358 26375
rect 7312 26226 7358 26272
rect 7312 26123 7358 26169
rect 7312 26019 7358 26065
rect 7556 26947 7602 26993
rect 7556 26844 7602 26890
rect 7556 26741 7602 26787
rect 7556 26638 7602 26684
rect 7556 26535 7602 26581
rect 7556 26432 7602 26478
rect 7556 26329 7602 26375
rect 7556 26226 7602 26272
rect 7556 26123 7602 26169
rect 7556 26019 7602 26065
rect 7800 26947 7846 26993
rect 7800 26844 7846 26890
rect 7800 26741 7846 26787
rect 7800 26638 7846 26684
rect 7800 26535 7846 26581
rect 7800 26432 7846 26478
rect 7800 26329 7846 26375
rect 7800 26226 7846 26272
rect 7800 26123 7846 26169
rect 7800 26019 7846 26065
rect 8044 26947 8090 26993
rect 8044 26844 8090 26890
rect 8044 26741 8090 26787
rect 8044 26638 8090 26684
rect 8044 26535 8090 26581
rect 8044 26432 8090 26478
rect 8044 26329 8090 26375
rect 8044 26226 8090 26272
rect 8044 26123 8090 26169
rect 8044 26019 8090 26065
<< mvpdiffc >>
rect 2590 28858 2636 28904
rect 2590 28755 2636 28801
rect 2590 28652 2636 28698
rect 2590 28549 2636 28595
rect 2590 28446 2636 28492
rect 2590 28343 2636 28389
rect 2590 28240 2636 28286
rect 2590 28137 2636 28183
rect 2590 28034 2636 28080
rect 2590 27930 2636 27976
rect 2834 28858 2880 28904
rect 2834 28755 2880 28801
rect 2834 28652 2880 28698
rect 2834 28549 2880 28595
rect 2834 28446 2880 28492
rect 2834 28343 2880 28389
rect 2834 28240 2880 28286
rect 2834 28137 2880 28183
rect 2834 28034 2880 28080
rect 2834 27930 2880 27976
rect 3078 28858 3124 28904
rect 3078 28755 3124 28801
rect 3078 28652 3124 28698
rect 3078 28549 3124 28595
rect 3078 28446 3124 28492
rect 3078 28343 3124 28389
rect 3078 28240 3124 28286
rect 3078 28137 3124 28183
rect 3078 28034 3124 28080
rect 3078 27930 3124 27976
rect 3322 28858 3368 28904
rect 3322 28755 3368 28801
rect 3322 28652 3368 28698
rect 3322 28549 3368 28595
rect 3322 28446 3368 28492
rect 3322 28343 3368 28389
rect 3322 28240 3368 28286
rect 3322 28137 3368 28183
rect 3322 28034 3368 28080
rect 3322 27930 3368 27976
rect 3566 28858 3612 28904
rect 3566 28755 3612 28801
rect 3566 28652 3612 28698
rect 3566 28549 3612 28595
rect 3566 28446 3612 28492
rect 3566 28343 3612 28389
rect 3566 28240 3612 28286
rect 3566 28137 3612 28183
rect 3566 28034 3612 28080
rect 3566 27930 3612 27976
rect 3810 28858 3856 28904
rect 3810 28755 3856 28801
rect 3810 28652 3856 28698
rect 3810 28549 3856 28595
rect 3810 28446 3856 28492
rect 3810 28343 3856 28389
rect 3810 28240 3856 28286
rect 3810 28137 3856 28183
rect 3810 28034 3856 28080
rect 3810 27930 3856 27976
rect 4054 28858 4100 28904
rect 4054 28755 4100 28801
rect 4054 28652 4100 28698
rect 4054 28549 4100 28595
rect 4054 28446 4100 28492
rect 4054 28343 4100 28389
rect 4054 28240 4100 28286
rect 4054 28137 4100 28183
rect 4054 28034 4100 28080
rect 4054 27930 4100 27976
rect 4298 28858 4344 28904
rect 4298 28755 4344 28801
rect 4298 28652 4344 28698
rect 4298 28549 4344 28595
rect 4298 28446 4344 28492
rect 4298 28343 4344 28389
rect 4298 28240 4344 28286
rect 4298 28137 4344 28183
rect 4298 28034 4344 28080
rect 4298 27930 4344 27976
rect 4470 28858 4516 28904
rect 4470 28755 4516 28801
rect 4470 28652 4516 28698
rect 4470 28549 4516 28595
rect 4470 28446 4516 28492
rect 4470 28343 4516 28389
rect 4470 28240 4516 28286
rect 4470 28137 4516 28183
rect 4470 28034 4516 28080
rect 4470 27930 4516 27976
rect 4714 28858 4760 28904
rect 4714 28755 4760 28801
rect 4714 28652 4760 28698
rect 4714 28549 4760 28595
rect 4714 28446 4760 28492
rect 4714 28343 4760 28389
rect 4714 28240 4760 28286
rect 4714 28137 4760 28183
rect 4714 28034 4760 28080
rect 4714 27930 4760 27976
rect 4958 28858 5004 28904
rect 4958 28755 5004 28801
rect 4958 28652 5004 28698
rect 4958 28549 5004 28595
rect 4958 28446 5004 28492
rect 4958 28343 5004 28389
rect 4958 28240 5004 28286
rect 4958 28137 5004 28183
rect 4958 28034 5004 28080
rect 4958 27930 5004 27976
rect 5202 28858 5248 28904
rect 5202 28755 5248 28801
rect 5202 28652 5248 28698
rect 5202 28549 5248 28595
rect 5202 28446 5248 28492
rect 5202 28343 5248 28389
rect 5202 28240 5248 28286
rect 5202 28137 5248 28183
rect 5202 28034 5248 28080
rect 5202 27930 5248 27976
rect 5446 28858 5492 28904
rect 5446 28755 5492 28801
rect 5446 28652 5492 28698
rect 5446 28549 5492 28595
rect 5446 28446 5492 28492
rect 5446 28343 5492 28389
rect 5446 28240 5492 28286
rect 5446 28137 5492 28183
rect 5446 28034 5492 28080
rect 5446 27930 5492 27976
rect 5690 28858 5736 28904
rect 5690 28755 5736 28801
rect 5690 28652 5736 28698
rect 5690 28549 5736 28595
rect 5690 28446 5736 28492
rect 5690 28343 5736 28389
rect 5690 28240 5736 28286
rect 5690 28137 5736 28183
rect 5690 28034 5736 28080
rect 5690 27930 5736 27976
rect 5934 28858 5980 28904
rect 5934 28755 5980 28801
rect 5934 28652 5980 28698
rect 5934 28549 5980 28595
rect 5934 28446 5980 28492
rect 5934 28343 5980 28389
rect 5934 28240 5980 28286
rect 5934 28137 5980 28183
rect 5934 28034 5980 28080
rect 5934 27930 5980 27976
rect 6178 28858 6224 28904
rect 6178 28755 6224 28801
rect 6178 28652 6224 28698
rect 6178 28549 6224 28595
rect 6178 28446 6224 28492
rect 6178 28343 6224 28389
rect 6178 28240 6224 28286
rect 6178 28137 6224 28183
rect 6178 28034 6224 28080
rect 6178 27930 6224 27976
rect 6422 28858 6468 28904
rect 6422 28755 6468 28801
rect 6422 28652 6468 28698
rect 6422 28549 6468 28595
rect 6422 28446 6468 28492
rect 6422 28343 6468 28389
rect 6422 28240 6468 28286
rect 6422 28137 6468 28183
rect 6422 28034 6468 28080
rect 6422 27930 6468 27976
rect 6666 28858 6712 28904
rect 6666 28755 6712 28801
rect 6666 28652 6712 28698
rect 6666 28549 6712 28595
rect 6666 28446 6712 28492
rect 6666 28343 6712 28389
rect 6666 28240 6712 28286
rect 6666 28137 6712 28183
rect 6666 28034 6712 28080
rect 6666 27930 6712 27976
rect 6910 28858 6956 28904
rect 6910 28755 6956 28801
rect 6910 28652 6956 28698
rect 6910 28549 6956 28595
rect 6910 28446 6956 28492
rect 6910 28343 6956 28389
rect 6910 28240 6956 28286
rect 6910 28137 6956 28183
rect 6910 28034 6956 28080
rect 6910 27930 6956 27976
rect 7154 28858 7200 28904
rect 7154 28755 7200 28801
rect 7154 28652 7200 28698
rect 7154 28549 7200 28595
rect 7154 28446 7200 28492
rect 7154 28343 7200 28389
rect 7154 28240 7200 28286
rect 7154 28137 7200 28183
rect 7154 28034 7200 28080
rect 7154 27930 7200 27976
rect 7398 28858 7444 28904
rect 7398 28755 7444 28801
rect 7398 28652 7444 28698
rect 7398 28549 7444 28595
rect 7398 28446 7444 28492
rect 7398 28343 7444 28389
rect 7398 28240 7444 28286
rect 7398 28137 7444 28183
rect 7398 28034 7444 28080
rect 7398 27930 7444 27976
rect 7642 28858 7688 28904
rect 7642 28755 7688 28801
rect 7642 28652 7688 28698
rect 7642 28549 7688 28595
rect 7642 28446 7688 28492
rect 7642 28343 7688 28389
rect 7642 28240 7688 28286
rect 7642 28137 7688 28183
rect 7642 28034 7688 28080
rect 7642 27930 7688 27976
rect 7886 28858 7932 28904
rect 7886 28755 7932 28801
rect 7886 28652 7932 28698
rect 7886 28549 7932 28595
rect 7886 28446 7932 28492
rect 7886 28343 7932 28389
rect 7886 28240 7932 28286
rect 7886 28137 7932 28183
rect 7886 28034 7932 28080
rect 7886 27930 7932 27976
rect 8130 28858 8176 28904
rect 8130 28755 8176 28801
rect 8130 28652 8176 28698
rect 8130 28549 8176 28595
rect 8130 28446 8176 28492
rect 8130 28343 8176 28389
rect 8130 28240 8176 28286
rect 8130 28137 8176 28183
rect 8130 28034 8176 28080
rect 8130 27930 8176 27976
rect 8374 28858 8420 28904
rect 8374 28755 8420 28801
rect 8374 28652 8420 28698
rect 8374 28549 8420 28595
rect 8374 28446 8420 28492
rect 8374 28343 8420 28389
rect 8374 28240 8420 28286
rect 8374 28137 8420 28183
rect 8374 28034 8420 28080
rect 8374 27930 8420 27976
rect 8618 28858 8664 28904
rect 8618 28755 8664 28801
rect 8618 28652 8664 28698
rect 8618 28549 8664 28595
rect 8618 28446 8664 28492
rect 8618 28343 8664 28389
rect 8618 28240 8664 28286
rect 8618 28137 8664 28183
rect 8618 28034 8664 28080
rect 8618 27930 8664 27976
rect 8862 28858 8908 28904
rect 8862 28755 8908 28801
rect 8862 28652 8908 28698
rect 8862 28549 8908 28595
rect 8862 28446 8908 28492
rect 8862 28343 8908 28389
rect 8862 28240 8908 28286
rect 8862 28137 8908 28183
rect 8862 28034 8908 28080
rect 8862 27930 8908 27976
rect 9106 28858 9152 28904
rect 9106 28755 9152 28801
rect 9106 28652 9152 28698
rect 9106 28549 9152 28595
rect 9106 28446 9152 28492
rect 9106 28343 9152 28389
rect 9106 28240 9152 28286
rect 9106 28137 9152 28183
rect 9106 28034 9152 28080
rect 9106 27930 9152 27976
rect 9350 28858 9396 28904
rect 9350 28755 9396 28801
rect 9350 28652 9396 28698
rect 9350 28549 9396 28595
rect 9350 28446 9396 28492
rect 9350 28343 9396 28389
rect 9350 28240 9396 28286
rect 9350 28137 9396 28183
rect 9350 28034 9396 28080
rect 9350 27930 9396 27976
rect 9594 28858 9640 28904
rect 9594 28755 9640 28801
rect 9594 28652 9640 28698
rect 9594 28549 9640 28595
rect 9594 28446 9640 28492
rect 9594 28343 9640 28389
rect 9594 28240 9640 28286
rect 9594 28137 9640 28183
rect 9594 28034 9640 28080
rect 9594 27930 9640 27976
rect 9838 28858 9884 28904
rect 9838 28755 9884 28801
rect 9838 28652 9884 28698
rect 9838 28549 9884 28595
rect 9838 28446 9884 28492
rect 9838 28343 9884 28389
rect 9838 28240 9884 28286
rect 9838 28137 9884 28183
rect 9838 28034 9884 28080
rect 9838 27930 9884 27976
rect 10082 28858 10128 28904
rect 10082 28755 10128 28801
rect 10082 28652 10128 28698
rect 10082 28549 10128 28595
rect 10082 28446 10128 28492
rect 10082 28343 10128 28389
rect 10082 28240 10128 28286
rect 10082 28137 10128 28183
rect 10082 28034 10128 28080
rect 10082 27930 10128 27976
rect 10326 28858 10372 28904
rect 10326 28755 10372 28801
rect 10326 28652 10372 28698
rect 10326 28549 10372 28595
rect 10326 28446 10372 28492
rect 10326 28343 10372 28389
rect 10326 28240 10372 28286
rect 10326 28137 10372 28183
rect 10326 28034 10372 28080
rect 10326 27930 10372 27976
<< psubdiff >>
rect 2253 27485 10709 27507
rect 2253 27439 3746 27485
rect 6518 27439 6887 27485
rect 10223 27439 10709 27485
rect 2253 27417 10709 27439
rect 2253 27156 2343 27417
rect 2253 25888 2275 27156
rect 2321 25888 2343 27156
rect 10619 27156 10709 27417
rect 2253 25802 2343 25888
rect 10619 25888 10641 27156
rect 10687 25888 10709 27156
rect 10619 25802 10709 25888
rect 2253 25780 10709 25802
rect 2253 25734 2275 25780
rect 6739 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10709 25780
rect 2253 25712 10709 25734
<< nsubdiff >>
rect 2253 29188 10709 29210
rect 2253 29142 2275 29188
rect 10687 29142 10709 29188
rect 2253 29120 10709 29142
rect 2253 29034 2343 29120
rect 2253 27860 2275 29034
rect 2321 27860 2343 29034
rect 10619 29034 10709 29120
rect 2253 27838 2343 27860
rect 10619 27860 10641 29034
rect 10687 27860 10709 29034
rect 10619 27838 10709 27860
<< psubdiffcont >>
rect 3746 27439 6518 27485
rect 6887 27439 10223 27485
rect 2275 25888 2321 27156
rect 10641 25888 10687 27156
rect 2275 25734 6739 25780
rect 6975 25734 7209 25780
rect 7445 25734 7679 25780
rect 8009 25734 10687 25780
<< nsubdiffcont >>
rect 2275 29142 10687 29188
rect 2275 27860 2321 29034
rect 10641 27860 10687 29034
<< polysilicon >>
rect 2665 28917 2805 28961
rect 2909 28917 3049 28961
rect 3153 28917 3293 28961
rect 3397 28917 3537 28961
rect 3641 28917 3781 28961
rect 3885 28917 4025 28961
rect 4129 28917 4269 28961
rect 4545 28917 4685 28961
rect 4789 28917 4929 28961
rect 5033 28917 5173 28961
rect 5277 28917 5417 28961
rect 5521 28917 5661 28961
rect 5765 28917 5905 28961
rect 6009 28917 6149 28961
rect 6253 28917 6393 28961
rect 6497 28917 6637 28961
rect 6741 28917 6881 28961
rect 6985 28917 7125 28961
rect 7229 28917 7369 28961
rect 7473 28917 7613 28961
rect 7717 28917 7857 28961
rect 7961 28917 8101 28961
rect 8205 28917 8345 28961
rect 8449 28917 8589 28961
rect 8693 28917 8833 28961
rect 8937 28917 9077 28961
rect 9181 28917 9321 28961
rect 9425 28917 9565 28961
rect 9669 28917 9809 28961
rect 9913 28917 10053 28961
rect 10157 28917 10297 28961
rect 2665 27729 2805 27917
rect 2909 27729 3049 27917
rect 3153 27729 3293 27917
rect 3397 27729 3537 27917
rect 2665 27710 3537 27729
rect 2665 27664 2749 27710
rect 3453 27664 3537 27710
rect 2665 27645 3537 27664
rect 3641 27729 3781 27917
rect 3885 27729 4025 27917
rect 4129 27729 4269 27917
rect 3641 27710 4269 27729
rect 3641 27664 3697 27710
rect 4213 27664 4269 27710
rect 3641 27645 4269 27664
rect 4545 27729 4685 27917
rect 4789 27729 4929 27917
rect 5033 27729 5173 27917
rect 5277 27729 5417 27917
rect 5521 27729 5661 27917
rect 5765 27729 5905 27917
rect 6009 27729 6149 27917
rect 6253 27729 6393 27917
rect 6497 27729 6637 27917
rect 6741 27729 6881 27917
rect 6985 27729 7125 27917
rect 7229 27729 7369 27917
rect 7473 27729 7613 27917
rect 7717 27729 7857 27917
rect 7961 27729 8101 27917
rect 8205 27729 8345 27917
rect 8449 27729 8589 27917
rect 8693 27729 8833 27917
rect 8937 27729 9077 27917
rect 9181 27729 9321 27917
rect 9425 27729 9565 27917
rect 9669 27729 9809 27917
rect 9913 27729 10053 27917
rect 10157 27729 10297 27917
rect 4545 27710 10297 27729
rect 4545 27664 4578 27710
rect 10264 27664 10297 27710
rect 4545 27645 10297 27664
rect 5191 27259 6551 27278
rect 5191 27213 5237 27259
rect 6505 27213 6551 27259
rect 5191 27194 6551 27213
rect 4053 27131 4269 27150
rect 4053 27085 4072 27131
rect 4212 27085 4269 27131
rect 4053 27066 4269 27085
rect 4129 27006 4269 27066
rect 5191 27006 5331 27194
rect 5435 27006 5575 27194
rect 5679 27006 5819 27194
rect 5923 27006 6063 27194
rect 6167 27006 6307 27194
rect 6411 27006 6551 27194
rect 6655 27259 8015 27278
rect 6655 27213 6701 27259
rect 7969 27213 8015 27259
rect 6655 27194 8015 27213
rect 6655 27006 6795 27194
rect 6899 27006 7039 27194
rect 7143 27006 7283 27194
rect 7387 27006 7527 27194
rect 7631 27006 7771 27194
rect 7875 27006 8015 27194
rect 4129 25962 4269 26006
rect 5191 25962 5331 26006
rect 5435 25962 5575 26006
rect 5679 25962 5819 26006
rect 5923 25962 6063 26006
rect 6167 25962 6307 26006
rect 6411 25962 6551 26006
rect 6655 25962 6795 26006
rect 6899 25962 7039 26006
rect 7143 25962 7283 26006
rect 7387 25962 7527 26006
rect 7631 25962 7771 26006
rect 7875 25962 8015 26006
<< polycontact >>
rect 2749 27664 3453 27710
rect 3697 27664 4213 27710
rect 4578 27664 10264 27710
rect 5237 27213 6505 27259
rect 4072 27085 4212 27131
rect 6701 27213 7969 27259
<< metal1 >>
rect -321 45914 -245 45926
rect -321 42118 -309 45914
rect -257 42118 -245 45914
rect -116 45914 1104 45926
rect -116 45862 -104 45914
rect 1092 45862 1104 45914
rect -116 45850 1104 45862
rect 1784 45914 3732 45926
rect 1784 45862 1796 45914
rect 3720 45862 3732 45914
rect 1784 45850 3732 45862
rect 4154 45914 6102 45926
rect 4154 45862 4166 45914
rect 6090 45862 6102 45914
rect 4154 45850 6102 45862
rect 6860 45914 8808 45926
rect 6860 45862 6872 45914
rect 8796 45862 8808 45914
rect 6860 45850 8808 45862
rect 9230 45914 11178 45926
rect 9230 45862 9242 45914
rect 11166 45862 11178 45914
rect 9230 45850 11178 45862
rect 11871 45914 13091 45926
rect 11871 45862 11883 45914
rect 13079 45862 13091 45914
rect 11871 45850 13091 45862
rect 13207 45914 13283 45926
rect -321 42106 -245 42118
rect 191 42174 1099 42186
rect 191 42122 203 42174
rect 1087 42122 1099 42174
rect 191 42110 1099 42122
rect 1784 42174 3732 42186
rect 1784 42122 1796 42174
rect 3720 42122 3732 42174
rect 1784 42110 3732 42122
rect 4154 42174 6102 42186
rect 4154 42122 4166 42174
rect 6090 42122 6102 42174
rect 4154 42110 6102 42122
rect 6860 42174 8808 42186
rect 6860 42122 6872 42174
rect 8796 42122 8808 42174
rect 6860 42110 8808 42122
rect 9230 42174 11178 42186
rect 9230 42122 9242 42174
rect 11166 42122 11178 42174
rect 9230 42110 11178 42122
rect 11871 42174 13091 42186
rect 11871 42122 11883 42174
rect 13079 42122 13091 42174
rect 11871 42110 13091 42122
rect 13207 42118 13219 45914
rect 13271 42118 13283 45914
rect 13207 42106 13283 42118
rect 1483 41733 1663 41745
rect 1483 41577 1495 41733
rect 1651 41577 1663 41733
rect 1483 41565 1663 41577
rect 3853 41733 4033 41745
rect 3853 41577 3865 41733
rect 4021 41577 4033 41733
rect 3853 41565 4033 41577
rect 6235 41733 6727 41745
rect 6235 41577 6247 41733
rect 6715 41577 6727 41733
rect 6235 41565 6727 41577
rect 8929 41733 9109 41745
rect 8929 41577 8941 41733
rect 9097 41577 9109 41733
rect 8929 41565 9109 41577
rect 11299 41733 11479 41745
rect 11299 41577 11311 41733
rect 11467 41577 11479 41733
rect 11299 41565 11479 41577
rect 1483 36000 1663 36012
rect 1483 35324 1495 36000
rect 1651 35324 1663 36000
rect 1483 35312 1663 35324
rect 3853 36000 4033 36012
rect 3853 35324 3865 36000
rect 4021 35324 4033 36000
rect 3853 35312 4033 35324
rect 6257 35998 6705 36010
rect 6257 35946 6269 35998
rect 6321 35946 6393 35998
rect 6445 35946 6517 35998
rect 6569 35946 6641 35998
rect 6693 35946 6705 35998
rect 6257 35874 6705 35946
rect 6257 35822 6269 35874
rect 6321 35822 6393 35874
rect 6445 35822 6517 35874
rect 6569 35822 6641 35874
rect 6693 35822 6705 35874
rect 6257 35750 6705 35822
rect 6257 35698 6269 35750
rect 6321 35698 6393 35750
rect 6445 35698 6517 35750
rect 6569 35698 6641 35750
rect 6693 35698 6705 35750
rect 6257 35626 6705 35698
rect 6257 35574 6269 35626
rect 6321 35574 6393 35626
rect 6445 35574 6517 35626
rect 6569 35574 6641 35626
rect 6693 35574 6705 35626
rect 6257 35502 6705 35574
rect 6257 35450 6269 35502
rect 6321 35450 6393 35502
rect 6445 35450 6517 35502
rect 6569 35450 6641 35502
rect 6693 35450 6705 35502
rect 6257 35378 6705 35450
rect 6257 35326 6269 35378
rect 6321 35326 6393 35378
rect 6445 35326 6517 35378
rect 6569 35326 6641 35378
rect 6693 35326 6705 35378
rect 6257 35314 6705 35326
rect 8929 36000 9109 36012
rect 8929 35324 8941 36000
rect 9097 35324 9109 36000
rect 8929 35312 9109 35324
rect 11299 36000 11479 36012
rect 11299 35324 11311 36000
rect 11467 35324 11479 36000
rect 11299 35312 11479 35324
rect -50 27721 110 30038
rect 1483 29649 1663 29661
rect 1483 29493 1495 29649
rect 1651 29493 1663 29649
rect 1483 29481 1663 29493
rect 3853 29649 4033 29661
rect 3853 29493 3865 29649
rect 4021 29493 4033 29649
rect 3853 29481 4033 29493
rect 6235 29649 6727 29661
rect 6235 29493 6247 29649
rect 6715 29493 6727 29649
rect 6235 29481 6727 29493
rect 8929 29649 9109 29661
rect 8929 29493 8941 29649
rect 9097 29493 9109 29649
rect 8929 29481 9109 29493
rect 11299 29649 11479 29661
rect 11299 29493 11311 29649
rect 11467 29493 11479 29649
rect 11299 29481 11479 29493
rect 2264 29188 10698 29199
rect 2264 29142 2275 29188
rect 10687 29142 10698 29188
rect 2264 29034 2276 29142
rect 2328 29131 10698 29142
rect 2264 27860 2275 29034
rect 2328 27861 2340 29131
rect 2575 29125 2651 29131
rect 2575 27929 2587 29125
rect 2639 27929 2651 29125
rect 3063 29125 3139 29131
rect 2575 27917 2651 27929
rect 2819 28904 2895 28917
rect 2819 28858 2834 28904
rect 2880 28858 2895 28904
rect 2819 28801 2895 28858
rect 2819 28755 2834 28801
rect 2880 28755 2895 28801
rect 2819 28698 2895 28755
rect 2819 28652 2834 28698
rect 2880 28652 2895 28698
rect 2819 28595 2895 28652
rect 2819 28549 2834 28595
rect 2880 28549 2895 28595
rect 2819 28492 2895 28549
rect 2819 28446 2834 28492
rect 2880 28446 2895 28492
rect 2819 28389 2895 28446
rect 2819 28343 2834 28389
rect 2880 28343 2895 28389
rect 2819 28286 2895 28343
rect 2819 28240 2834 28286
rect 2880 28240 2895 28286
rect 2819 28183 2895 28240
rect 2819 28137 2834 28183
rect 2880 28137 2895 28183
rect 2819 28080 2895 28137
rect 2819 28034 2834 28080
rect 2880 28034 2895 28080
rect 2819 27976 2895 28034
rect 2819 27930 2834 27976
rect 2880 27930 2895 27976
rect 2321 27860 2340 27861
rect 2264 27849 2340 27860
rect 2819 27857 2895 27930
rect 3063 27929 3075 29125
rect 3127 27929 3139 29125
rect 3551 29125 3627 29131
rect 3063 27917 3139 27929
rect 3307 28904 3383 28917
rect 3307 28858 3322 28904
rect 3368 28858 3383 28904
rect 3307 28801 3383 28858
rect 3307 28755 3322 28801
rect 3368 28755 3383 28801
rect 3307 28698 3383 28755
rect 3307 28652 3322 28698
rect 3368 28652 3383 28698
rect 3307 28595 3383 28652
rect 3307 28549 3322 28595
rect 3368 28549 3383 28595
rect 3307 28492 3383 28549
rect 3307 28446 3322 28492
rect 3368 28446 3383 28492
rect 3307 28389 3383 28446
rect 3307 28343 3322 28389
rect 3368 28343 3383 28389
rect 3307 28286 3383 28343
rect 3307 28240 3322 28286
rect 3368 28240 3383 28286
rect 3307 28183 3383 28240
rect 3307 28137 3322 28183
rect 3368 28137 3383 28183
rect 3307 28080 3383 28137
rect 3307 28034 3322 28080
rect 3368 28034 3383 28080
rect 3307 27976 3383 28034
rect 3307 27930 3322 27976
rect 3368 27930 3383 27976
rect 3307 27857 3383 27930
rect 3551 27929 3563 29125
rect 3615 27929 3627 29125
rect 3551 27917 3627 27929
rect 3795 28904 3871 28917
rect 3795 28858 3810 28904
rect 3856 28858 3871 28904
rect 3795 28801 3871 28858
rect 3795 28755 3810 28801
rect 3856 28755 3871 28801
rect 3795 28698 3871 28755
rect 3795 28652 3810 28698
rect 3856 28652 3871 28698
rect 3795 28595 3871 28652
rect 3795 28549 3810 28595
rect 3856 28549 3871 28595
rect 3795 28492 3871 28549
rect 3795 28446 3810 28492
rect 3856 28446 3871 28492
rect 3795 28389 3871 28446
rect 3795 28343 3810 28389
rect 3856 28343 3871 28389
rect 3795 28286 3871 28343
rect 3795 28240 3810 28286
rect 3856 28240 3871 28286
rect 3795 28183 3871 28240
rect 3795 28137 3810 28183
rect 3856 28137 3871 28183
rect 3795 28080 3871 28137
rect 3795 28034 3810 28080
rect 3856 28034 3871 28080
rect 3795 27976 3871 28034
rect 3795 27930 3810 27976
rect 3856 27930 3871 27976
rect 3795 27857 3871 27930
rect 4039 28904 4115 29131
rect 4455 29125 4531 29131
rect 4039 28858 4054 28904
rect 4100 28858 4115 28904
rect 4039 28801 4115 28858
rect 4039 28755 4054 28801
rect 4100 28755 4115 28801
rect 4039 28698 4115 28755
rect 4039 28652 4054 28698
rect 4100 28652 4115 28698
rect 4039 28595 4115 28652
rect 4039 28549 4054 28595
rect 4100 28549 4115 28595
rect 4039 28492 4115 28549
rect 4039 28446 4054 28492
rect 4100 28446 4115 28492
rect 4039 28389 4115 28446
rect 4039 28343 4054 28389
rect 4100 28343 4115 28389
rect 4039 28286 4115 28343
rect 4039 28240 4054 28286
rect 4100 28240 4115 28286
rect 4039 28183 4115 28240
rect 4039 28137 4054 28183
rect 4100 28137 4115 28183
rect 4039 28080 4115 28137
rect 4039 28034 4054 28080
rect 4100 28034 4115 28080
rect 4039 27976 4115 28034
rect 4039 27930 4054 27976
rect 4100 27930 4115 27976
rect 4039 27917 4115 27930
rect 4283 28904 4359 28917
rect 4283 28858 4298 28904
rect 4344 28858 4359 28904
rect 4283 28801 4359 28858
rect 4283 28755 4298 28801
rect 4344 28755 4359 28801
rect 4283 28698 4359 28755
rect 4283 28652 4298 28698
rect 4344 28652 4359 28698
rect 4283 28595 4359 28652
rect 4283 28549 4298 28595
rect 4344 28549 4359 28595
rect 4283 28492 4359 28549
rect 4283 28446 4298 28492
rect 4344 28446 4359 28492
rect 4283 28389 4359 28446
rect 4283 28343 4298 28389
rect 4344 28343 4359 28389
rect 4283 28286 4359 28343
rect 4283 28240 4298 28286
rect 4344 28240 4359 28286
rect 4283 28183 4359 28240
rect 4283 28137 4298 28183
rect 4344 28137 4359 28183
rect 4283 28080 4359 28137
rect 4283 28034 4298 28080
rect 4344 28034 4359 28080
rect 4283 27976 4359 28034
rect 4283 27930 4298 27976
rect 4344 27930 4359 27976
rect 4283 27857 4359 27930
rect 4455 27929 4467 29125
rect 4519 27929 4531 29125
rect 4943 29125 5019 29131
rect 4455 27917 4531 27929
rect 4699 28904 4775 28917
rect 4699 28858 4714 28904
rect 4760 28858 4775 28904
rect 4699 28801 4775 28858
rect 4699 28755 4714 28801
rect 4760 28755 4775 28801
rect 4699 28698 4775 28755
rect 4699 28652 4714 28698
rect 4760 28652 4775 28698
rect 4699 28595 4775 28652
rect 4699 28549 4714 28595
rect 4760 28549 4775 28595
rect 4699 28492 4775 28549
rect 4699 28446 4714 28492
rect 4760 28446 4775 28492
rect 4699 28389 4775 28446
rect 4699 28343 4714 28389
rect 4760 28343 4775 28389
rect 4699 28286 4775 28343
rect 4699 28240 4714 28286
rect 4760 28240 4775 28286
rect 4699 28183 4775 28240
rect 4699 28137 4714 28183
rect 4760 28137 4775 28183
rect 4699 28080 4775 28137
rect 4699 28034 4714 28080
rect 4760 28034 4775 28080
rect 4699 27976 4775 28034
rect 4699 27930 4714 27976
rect 4760 27930 4775 27976
rect 2819 27781 3627 27857
rect 3795 27781 4359 27857
rect 4699 27857 4775 27930
rect 4943 27929 4955 29125
rect 5007 27929 5019 29125
rect 5431 29125 5507 29131
rect 4943 27917 5019 27929
rect 5187 28904 5263 28917
rect 5187 28858 5202 28904
rect 5248 28858 5263 28904
rect 5187 28801 5263 28858
rect 5187 28755 5202 28801
rect 5248 28755 5263 28801
rect 5187 28698 5263 28755
rect 5187 28652 5202 28698
rect 5248 28652 5263 28698
rect 5187 28595 5263 28652
rect 5187 28549 5202 28595
rect 5248 28549 5263 28595
rect 5187 28492 5263 28549
rect 5187 28446 5202 28492
rect 5248 28446 5263 28492
rect 5187 28389 5263 28446
rect 5187 28343 5202 28389
rect 5248 28343 5263 28389
rect 5187 28286 5263 28343
rect 5187 28240 5202 28286
rect 5248 28240 5263 28286
rect 5187 28183 5263 28240
rect 5187 28137 5202 28183
rect 5248 28137 5263 28183
rect 5187 28080 5263 28137
rect 5187 28034 5202 28080
rect 5248 28034 5263 28080
rect 5187 27976 5263 28034
rect 5187 27930 5202 27976
rect 5248 27930 5263 27976
rect 5187 27857 5263 27930
rect 5431 27929 5443 29125
rect 5495 27929 5507 29125
rect 5919 29125 5995 29131
rect 5431 27917 5507 27929
rect 5675 28904 5751 28917
rect 5675 28858 5690 28904
rect 5736 28858 5751 28904
rect 5675 28801 5751 28858
rect 5675 28755 5690 28801
rect 5736 28755 5751 28801
rect 5675 28698 5751 28755
rect 5675 28652 5690 28698
rect 5736 28652 5751 28698
rect 5675 28595 5751 28652
rect 5675 28549 5690 28595
rect 5736 28549 5751 28595
rect 5675 28492 5751 28549
rect 5675 28446 5690 28492
rect 5736 28446 5751 28492
rect 5675 28389 5751 28446
rect 5675 28343 5690 28389
rect 5736 28343 5751 28389
rect 5675 28286 5751 28343
rect 5675 28240 5690 28286
rect 5736 28240 5751 28286
rect 5675 28183 5751 28240
rect 5675 28137 5690 28183
rect 5736 28137 5751 28183
rect 5675 28080 5751 28137
rect 5675 28034 5690 28080
rect 5736 28034 5751 28080
rect 5675 27976 5751 28034
rect 5675 27930 5690 27976
rect 5736 27930 5751 27976
rect 5675 27857 5751 27930
rect 5919 27929 5931 29125
rect 5983 27929 5995 29125
rect 5919 27917 5995 27929
rect 6163 28904 6239 28917
rect 6163 28858 6178 28904
rect 6224 28858 6239 28904
rect 6163 28801 6239 28858
rect 6163 28755 6178 28801
rect 6224 28755 6239 28801
rect 6163 28698 6239 28755
rect 6163 28652 6178 28698
rect 6224 28652 6239 28698
rect 6163 28595 6239 28652
rect 6163 28549 6178 28595
rect 6224 28549 6239 28595
rect 6163 28492 6239 28549
rect 6163 28446 6178 28492
rect 6224 28446 6239 28492
rect 6163 28389 6239 28446
rect 6163 28343 6178 28389
rect 6224 28343 6239 28389
rect 6163 28286 6239 28343
rect 6163 28240 6178 28286
rect 6224 28240 6239 28286
rect 6163 28183 6239 28240
rect 6163 28137 6178 28183
rect 6224 28137 6239 28183
rect 6163 28080 6239 28137
rect 6163 28034 6178 28080
rect 6224 28034 6239 28080
rect 6163 27976 6239 28034
rect 6163 27930 6178 27976
rect 6224 27930 6239 27976
rect 6163 27857 6239 27930
rect 6407 28904 6483 29131
rect 6895 29125 6971 29131
rect 6407 28858 6422 28904
rect 6468 28858 6483 28904
rect 6407 28801 6483 28858
rect 6407 28755 6422 28801
rect 6468 28755 6483 28801
rect 6407 28698 6483 28755
rect 6407 28652 6422 28698
rect 6468 28652 6483 28698
rect 6407 28595 6483 28652
rect 6407 28549 6422 28595
rect 6468 28549 6483 28595
rect 6407 28492 6483 28549
rect 6407 28446 6422 28492
rect 6468 28446 6483 28492
rect 6407 28389 6483 28446
rect 6407 28343 6422 28389
rect 6468 28343 6483 28389
rect 6407 28286 6483 28343
rect 6407 28240 6422 28286
rect 6468 28240 6483 28286
rect 6407 28183 6483 28240
rect 6407 28137 6422 28183
rect 6468 28137 6483 28183
rect 6407 28080 6483 28137
rect 6407 28034 6422 28080
rect 6468 28034 6483 28080
rect 6407 27976 6483 28034
rect 6407 27930 6422 27976
rect 6468 27930 6483 27976
rect 6407 27917 6483 27930
rect 6651 28904 6727 28917
rect 6651 28858 6666 28904
rect 6712 28858 6727 28904
rect 6651 28801 6727 28858
rect 6651 28755 6666 28801
rect 6712 28755 6727 28801
rect 6651 28698 6727 28755
rect 6651 28652 6666 28698
rect 6712 28652 6727 28698
rect 6651 28595 6727 28652
rect 6651 28549 6666 28595
rect 6712 28549 6727 28595
rect 6651 28492 6727 28549
rect 6651 28446 6666 28492
rect 6712 28446 6727 28492
rect 6651 28389 6727 28446
rect 6651 28343 6666 28389
rect 6712 28343 6727 28389
rect 6651 28286 6727 28343
rect 6651 28240 6666 28286
rect 6712 28240 6727 28286
rect 6651 28183 6727 28240
rect 6651 28137 6666 28183
rect 6712 28137 6727 28183
rect 6651 28080 6727 28137
rect 6651 28034 6666 28080
rect 6712 28034 6727 28080
rect 6651 27976 6727 28034
rect 6651 27930 6666 27976
rect 6712 27930 6727 27976
rect 6651 27857 6727 27930
rect 6895 27929 6907 29125
rect 6959 27929 6971 29125
rect 7383 29125 7459 29131
rect 6895 27917 6971 27929
rect 7139 28904 7215 28917
rect 7139 28858 7154 28904
rect 7200 28858 7215 28904
rect 7139 28801 7215 28858
rect 7139 28755 7154 28801
rect 7200 28755 7215 28801
rect 7139 28698 7215 28755
rect 7139 28652 7154 28698
rect 7200 28652 7215 28698
rect 7139 28595 7215 28652
rect 7139 28549 7154 28595
rect 7200 28549 7215 28595
rect 7139 28492 7215 28549
rect 7139 28446 7154 28492
rect 7200 28446 7215 28492
rect 7139 28389 7215 28446
rect 7139 28343 7154 28389
rect 7200 28343 7215 28389
rect 7139 28286 7215 28343
rect 7139 28240 7154 28286
rect 7200 28240 7215 28286
rect 7139 28183 7215 28240
rect 7139 28137 7154 28183
rect 7200 28137 7215 28183
rect 7139 28080 7215 28137
rect 7139 28034 7154 28080
rect 7200 28034 7215 28080
rect 7139 27976 7215 28034
rect 7139 27930 7154 27976
rect 7200 27930 7215 27976
rect 7139 27857 7215 27930
rect 7383 27929 7395 29125
rect 7447 27929 7459 29125
rect 7871 29125 7947 29131
rect 7383 27917 7459 27929
rect 7627 28904 7703 28917
rect 7627 28858 7642 28904
rect 7688 28858 7703 28904
rect 7627 28801 7703 28858
rect 7627 28755 7642 28801
rect 7688 28755 7703 28801
rect 7627 28698 7703 28755
rect 7627 28652 7642 28698
rect 7688 28652 7703 28698
rect 7627 28595 7703 28652
rect 7627 28549 7642 28595
rect 7688 28549 7703 28595
rect 7627 28492 7703 28549
rect 7627 28446 7642 28492
rect 7688 28446 7703 28492
rect 7627 28389 7703 28446
rect 7627 28343 7642 28389
rect 7688 28343 7703 28389
rect 7627 28286 7703 28343
rect 7627 28240 7642 28286
rect 7688 28240 7703 28286
rect 7627 28183 7703 28240
rect 7627 28137 7642 28183
rect 7688 28137 7703 28183
rect 7627 28080 7703 28137
rect 7627 28034 7642 28080
rect 7688 28034 7703 28080
rect 7627 27976 7703 28034
rect 7627 27930 7642 27976
rect 7688 27930 7703 27976
rect 7627 27857 7703 27930
rect 7871 27929 7883 29125
rect 7935 27929 7947 29125
rect 8359 29125 8435 29131
rect 7871 27917 7947 27929
rect 8115 28904 8191 28917
rect 8115 28858 8130 28904
rect 8176 28858 8191 28904
rect 8115 28801 8191 28858
rect 8115 28755 8130 28801
rect 8176 28755 8191 28801
rect 8115 28698 8191 28755
rect 8115 28652 8130 28698
rect 8176 28652 8191 28698
rect 8115 28595 8191 28652
rect 8115 28549 8130 28595
rect 8176 28549 8191 28595
rect 8115 28492 8191 28549
rect 8115 28446 8130 28492
rect 8176 28446 8191 28492
rect 8115 28389 8191 28446
rect 8115 28343 8130 28389
rect 8176 28343 8191 28389
rect 8115 28286 8191 28343
rect 8115 28240 8130 28286
rect 8176 28240 8191 28286
rect 8115 28183 8191 28240
rect 8115 28137 8130 28183
rect 8176 28137 8191 28183
rect 8115 28080 8191 28137
rect 8115 28034 8130 28080
rect 8176 28034 8191 28080
rect 8115 27976 8191 28034
rect 8115 27930 8130 27976
rect 8176 27930 8191 27976
rect 8115 27857 8191 27930
rect 8359 27929 8371 29125
rect 8423 27929 8435 29125
rect 8359 27917 8435 27929
rect 8603 28904 8679 28917
rect 8603 28858 8618 28904
rect 8664 28858 8679 28904
rect 8603 28801 8679 28858
rect 8603 28755 8618 28801
rect 8664 28755 8679 28801
rect 8603 28698 8679 28755
rect 8603 28652 8618 28698
rect 8664 28652 8679 28698
rect 8603 28595 8679 28652
rect 8603 28549 8618 28595
rect 8664 28549 8679 28595
rect 8603 28492 8679 28549
rect 8603 28446 8618 28492
rect 8664 28446 8679 28492
rect 8603 28389 8679 28446
rect 8603 28343 8618 28389
rect 8664 28343 8679 28389
rect 8603 28286 8679 28343
rect 8603 28240 8618 28286
rect 8664 28240 8679 28286
rect 8603 28183 8679 28240
rect 8603 28137 8618 28183
rect 8664 28137 8679 28183
rect 8603 28080 8679 28137
rect 8603 28034 8618 28080
rect 8664 28034 8679 28080
rect 8603 27976 8679 28034
rect 8603 27930 8618 27976
rect 8664 27930 8679 27976
rect 8603 27857 8679 27930
rect 8847 28904 8923 29131
rect 9335 29125 9411 29131
rect 8847 28858 8862 28904
rect 8908 28858 8923 28904
rect 8847 28801 8923 28858
rect 8847 28755 8862 28801
rect 8908 28755 8923 28801
rect 8847 28698 8923 28755
rect 8847 28652 8862 28698
rect 8908 28652 8923 28698
rect 8847 28595 8923 28652
rect 8847 28549 8862 28595
rect 8908 28549 8923 28595
rect 8847 28492 8923 28549
rect 8847 28446 8862 28492
rect 8908 28446 8923 28492
rect 8847 28389 8923 28446
rect 8847 28343 8862 28389
rect 8908 28343 8923 28389
rect 8847 28286 8923 28343
rect 8847 28240 8862 28286
rect 8908 28240 8923 28286
rect 8847 28183 8923 28240
rect 8847 28137 8862 28183
rect 8908 28137 8923 28183
rect 8847 28080 8923 28137
rect 8847 28034 8862 28080
rect 8908 28034 8923 28080
rect 8847 27976 8923 28034
rect 8847 27930 8862 27976
rect 8908 27930 8923 27976
rect 8847 27917 8923 27930
rect 9091 28904 9167 28917
rect 9091 28858 9106 28904
rect 9152 28858 9167 28904
rect 9091 28801 9167 28858
rect 9091 28755 9106 28801
rect 9152 28755 9167 28801
rect 9091 28698 9167 28755
rect 9091 28652 9106 28698
rect 9152 28652 9167 28698
rect 9091 28595 9167 28652
rect 9091 28549 9106 28595
rect 9152 28549 9167 28595
rect 9091 28492 9167 28549
rect 9091 28446 9106 28492
rect 9152 28446 9167 28492
rect 9091 28389 9167 28446
rect 9091 28343 9106 28389
rect 9152 28343 9167 28389
rect 9091 28286 9167 28343
rect 9091 28240 9106 28286
rect 9152 28240 9167 28286
rect 9091 28183 9167 28240
rect 9091 28137 9106 28183
rect 9152 28137 9167 28183
rect 9091 28080 9167 28137
rect 9091 28034 9106 28080
rect 9152 28034 9167 28080
rect 9091 27976 9167 28034
rect 9091 27930 9106 27976
rect 9152 27930 9167 27976
rect 9091 27857 9167 27930
rect 9335 27929 9347 29125
rect 9399 27929 9411 29125
rect 9823 29125 9899 29131
rect 9335 27917 9411 27929
rect 9579 28904 9655 28917
rect 9579 28858 9594 28904
rect 9640 28858 9655 28904
rect 9579 28801 9655 28858
rect 9579 28755 9594 28801
rect 9640 28755 9655 28801
rect 9579 28698 9655 28755
rect 9579 28652 9594 28698
rect 9640 28652 9655 28698
rect 9579 28595 9655 28652
rect 9579 28549 9594 28595
rect 9640 28549 9655 28595
rect 9579 28492 9655 28549
rect 9579 28446 9594 28492
rect 9640 28446 9655 28492
rect 9579 28389 9655 28446
rect 9579 28343 9594 28389
rect 9640 28343 9655 28389
rect 9579 28286 9655 28343
rect 9579 28240 9594 28286
rect 9640 28240 9655 28286
rect 9579 28183 9655 28240
rect 9579 28137 9594 28183
rect 9640 28137 9655 28183
rect 9579 28080 9655 28137
rect 9579 28034 9594 28080
rect 9640 28034 9655 28080
rect 9579 27976 9655 28034
rect 9579 27930 9594 27976
rect 9640 27930 9655 27976
rect 9579 27857 9655 27930
rect 9823 27929 9835 29125
rect 9887 27929 9899 29125
rect 10311 29125 10387 29131
rect 9823 27917 9899 27929
rect 10067 28904 10143 28917
rect 10067 28858 10082 28904
rect 10128 28858 10143 28904
rect 10067 28801 10143 28858
rect 10067 28755 10082 28801
rect 10128 28755 10143 28801
rect 10067 28698 10143 28755
rect 10067 28652 10082 28698
rect 10128 28652 10143 28698
rect 10067 28595 10143 28652
rect 10067 28549 10082 28595
rect 10128 28549 10143 28595
rect 10067 28492 10143 28549
rect 10067 28446 10082 28492
rect 10128 28446 10143 28492
rect 10067 28389 10143 28446
rect 10067 28343 10082 28389
rect 10128 28343 10143 28389
rect 10067 28286 10143 28343
rect 10067 28240 10082 28286
rect 10128 28240 10143 28286
rect 10067 28183 10143 28240
rect 10067 28137 10082 28183
rect 10128 28137 10143 28183
rect 10067 28080 10143 28137
rect 10067 28034 10082 28080
rect 10128 28034 10143 28080
rect 10067 27976 10143 28034
rect 10067 27930 10082 27976
rect 10128 27930 10143 27976
rect 10067 27857 10143 27930
rect 10311 27929 10323 29125
rect 10375 27929 10387 29125
rect 10311 27917 10387 27929
rect 10622 29125 10698 29131
rect 10622 27929 10634 29125
rect 10686 29034 10698 29125
rect 10622 27917 10641 27929
rect 10630 27860 10641 27917
rect 10687 27860 10698 29034
rect 4699 27781 10433 27857
rect 10630 27849 10698 27860
rect 3551 27725 3627 27781
rect -50 27710 3464 27721
rect -50 27664 2749 27710
rect 3453 27664 3464 27710
rect -50 27521 3464 27664
rect 2264 27156 2332 27167
rect 2264 25888 2275 27156
rect 2321 25888 2332 27156
rect 3388 27146 3464 27521
rect 3551 27710 4224 27725
rect 3551 27664 3697 27710
rect 4213 27664 4224 27710
rect 3551 27649 4224 27664
rect 4283 27721 4359 27781
rect 4283 27710 10275 27721
rect 4283 27664 4578 27710
rect 10264 27664 10275 27710
rect 3551 27274 3627 27649
rect 4283 27645 10275 27664
rect 3735 27485 6529 27496
rect 3735 27439 3746 27485
rect 6518 27439 6529 27485
rect 3735 27432 3865 27439
rect 4021 27432 6257 27439
rect 6517 27432 6529 27439
rect 3735 27428 6529 27432
rect 3853 27420 4033 27428
rect 6245 27420 6529 27428
rect 3551 27259 6516 27274
rect 3551 27213 5237 27259
rect 6505 27213 6516 27259
rect 3551 27198 6516 27213
rect 6652 27270 6728 27645
rect 6876 27485 10234 27496
rect 6876 27439 6887 27485
rect 10223 27439 10234 27485
rect 6876 27432 8941 27439
rect 9097 27432 10234 27439
rect 6876 27428 10234 27432
rect 8929 27420 9109 27428
rect 6652 27259 7980 27270
rect 6652 27213 6701 27259
rect 7969 27213 7980 27259
rect 6652 27202 7980 27213
rect 3388 27131 4223 27146
rect 3388 27085 4072 27131
rect 4212 27085 4223 27131
rect 3388 27070 4223 27085
rect 2264 25799 2332 25888
rect 4039 26993 4115 27006
rect 4039 26947 4054 26993
rect 4100 26947 4115 26993
rect 4039 26890 4115 26947
rect 4039 26844 4054 26890
rect 4100 26844 4115 26890
rect 4039 26787 4115 26844
rect 4039 26741 4054 26787
rect 4100 26741 4115 26787
rect 4039 26684 4115 26741
rect 4039 26638 4054 26684
rect 4100 26638 4115 26684
rect 4039 26581 4115 26638
rect 4039 26535 4054 26581
rect 4100 26535 4115 26581
rect 4039 26478 4115 26535
rect 4039 26432 4054 26478
rect 4100 26432 4115 26478
rect 4039 26375 4115 26432
rect 4039 26329 4054 26375
rect 4100 26329 4115 26375
rect 4039 26272 4115 26329
rect 4039 26226 4054 26272
rect 4100 26226 4115 26272
rect 4039 26169 4115 26226
rect 4039 26123 4054 26169
rect 4100 26123 4115 26169
rect 4039 26065 4115 26123
rect 4039 26019 4054 26065
rect 4100 26019 4115 26065
rect 4039 25799 4115 26019
rect 4283 26993 4359 27198
rect 6652 27142 6728 27202
rect 10357 27142 10433 27781
rect 5345 27066 6728 27142
rect 6809 27066 10433 27142
rect 10630 27156 10698 27167
rect 4283 26947 4298 26993
rect 4344 26947 4359 26993
rect 4283 26890 4359 26947
rect 4283 26844 4298 26890
rect 4344 26844 4359 26890
rect 4283 26787 4359 26844
rect 4283 26741 4298 26787
rect 4344 26741 4359 26787
rect 4283 26684 4359 26741
rect 4283 26638 4298 26684
rect 4344 26638 4359 26684
rect 4283 26581 4359 26638
rect 4283 26535 4298 26581
rect 4344 26535 4359 26581
rect 4283 26478 4359 26535
rect 4283 26432 4298 26478
rect 4344 26432 4359 26478
rect 4283 26375 4359 26432
rect 4283 26329 4298 26375
rect 4344 26329 4359 26375
rect 4283 26272 4359 26329
rect 4283 26226 4298 26272
rect 4344 26226 4359 26272
rect 4283 26169 4359 26226
rect 4283 26123 4298 26169
rect 4344 26123 4359 26169
rect 4283 26065 4359 26123
rect 4283 26019 4298 26065
rect 4344 26019 4359 26065
rect 4283 26006 4359 26019
rect 5101 26993 5177 27006
rect 5101 26947 5116 26993
rect 5162 26947 5177 26993
rect 5101 26890 5177 26947
rect 5101 26844 5116 26890
rect 5162 26844 5177 26890
rect 5101 26787 5177 26844
rect 5101 26741 5116 26787
rect 5162 26741 5177 26787
rect 5101 26684 5177 26741
rect 5101 26638 5116 26684
rect 5162 26638 5177 26684
rect 5101 26581 5177 26638
rect 5101 26535 5116 26581
rect 5162 26535 5177 26581
rect 5101 26478 5177 26535
rect 5101 26432 5116 26478
rect 5162 26432 5177 26478
rect 5101 26375 5177 26432
rect 5101 26329 5116 26375
rect 5162 26329 5177 26375
rect 5101 26272 5177 26329
rect 5101 26226 5116 26272
rect 5162 26226 5177 26272
rect 5101 26169 5177 26226
rect 5101 26123 5116 26169
rect 5162 26123 5177 26169
rect 5101 26065 5177 26123
rect 5101 26019 5116 26065
rect 5162 26019 5177 26065
rect 1473 25791 2332 25799
rect 3853 25791 4115 25799
rect 5101 25791 5177 26019
rect 5345 26993 5421 27066
rect 5345 26947 5360 26993
rect 5406 26947 5421 26993
rect 5345 26890 5421 26947
rect 5345 26844 5360 26890
rect 5406 26844 5421 26890
rect 5345 26787 5421 26844
rect 5345 26741 5360 26787
rect 5406 26741 5421 26787
rect 5345 26684 5421 26741
rect 5345 26638 5360 26684
rect 5406 26638 5421 26684
rect 5345 26581 5421 26638
rect 5345 26535 5360 26581
rect 5406 26535 5421 26581
rect 5345 26478 5421 26535
rect 5345 26432 5360 26478
rect 5406 26432 5421 26478
rect 5345 26375 5421 26432
rect 5345 26329 5360 26375
rect 5406 26329 5421 26375
rect 5345 26272 5421 26329
rect 5345 26226 5360 26272
rect 5406 26226 5421 26272
rect 5345 26169 5421 26226
rect 5345 26123 5360 26169
rect 5406 26123 5421 26169
rect 5345 26065 5421 26123
rect 5345 26019 5360 26065
rect 5406 26019 5421 26065
rect 5345 26006 5421 26019
rect 5589 26993 5665 27006
rect 5589 26947 5604 26993
rect 5650 26947 5665 26993
rect 5589 26890 5665 26947
rect 5589 26844 5604 26890
rect 5650 26844 5665 26890
rect 5589 26787 5665 26844
rect 5589 26741 5604 26787
rect 5650 26741 5665 26787
rect 5589 26684 5665 26741
rect 5589 26638 5604 26684
rect 5650 26638 5665 26684
rect 5589 26581 5665 26638
rect 5589 26535 5604 26581
rect 5650 26535 5665 26581
rect 5589 26478 5665 26535
rect 5589 26432 5604 26478
rect 5650 26432 5665 26478
rect 5589 26375 5665 26432
rect 5589 26329 5604 26375
rect 5650 26329 5665 26375
rect 5589 26272 5665 26329
rect 5589 26226 5604 26272
rect 5650 26226 5665 26272
rect 5589 26169 5665 26226
rect 5589 26123 5604 26169
rect 5650 26123 5665 26169
rect 5589 26065 5665 26123
rect 5589 26019 5604 26065
rect 5650 26019 5665 26065
rect 5589 25791 5665 26019
rect 5833 26993 5909 27066
rect 5833 26947 5848 26993
rect 5894 26947 5909 26993
rect 5833 26890 5909 26947
rect 5833 26844 5848 26890
rect 5894 26844 5909 26890
rect 5833 26787 5909 26844
rect 5833 26741 5848 26787
rect 5894 26741 5909 26787
rect 5833 26684 5909 26741
rect 5833 26638 5848 26684
rect 5894 26638 5909 26684
rect 5833 26581 5909 26638
rect 5833 26535 5848 26581
rect 5894 26535 5909 26581
rect 5833 26478 5909 26535
rect 5833 26432 5848 26478
rect 5894 26432 5909 26478
rect 5833 26375 5909 26432
rect 5833 26329 5848 26375
rect 5894 26329 5909 26375
rect 5833 26272 5909 26329
rect 5833 26226 5848 26272
rect 5894 26226 5909 26272
rect 5833 26169 5909 26226
rect 5833 26123 5848 26169
rect 5894 26123 5909 26169
rect 5833 26065 5909 26123
rect 5833 26019 5848 26065
rect 5894 26019 5909 26065
rect 5833 26006 5909 26019
rect 6077 26993 6153 27006
rect 6077 26947 6092 26993
rect 6138 26947 6153 26993
rect 6077 26890 6153 26947
rect 6077 26844 6092 26890
rect 6138 26844 6153 26890
rect 6077 26787 6153 26844
rect 6077 26741 6092 26787
rect 6138 26741 6153 26787
rect 6077 26684 6153 26741
rect 6077 26638 6092 26684
rect 6138 26638 6153 26684
rect 6077 26581 6153 26638
rect 6077 26535 6092 26581
rect 6138 26535 6153 26581
rect 6077 26478 6153 26535
rect 6077 26432 6092 26478
rect 6138 26432 6153 26478
rect 6077 26375 6153 26432
rect 6077 26329 6092 26375
rect 6138 26329 6153 26375
rect 6077 26272 6153 26329
rect 6077 26226 6092 26272
rect 6138 26226 6153 26272
rect 6077 26169 6153 26226
rect 6077 26123 6092 26169
rect 6138 26123 6153 26169
rect 6077 26065 6153 26123
rect 6077 26019 6092 26065
rect 6138 26019 6153 26065
rect 6077 25791 6153 26019
rect 6321 26993 6397 27066
rect 6321 26947 6336 26993
rect 6382 26947 6397 26993
rect 6321 26890 6397 26947
rect 6321 26844 6336 26890
rect 6382 26844 6397 26890
rect 6321 26787 6397 26844
rect 6321 26741 6336 26787
rect 6382 26741 6397 26787
rect 6321 26684 6397 26741
rect 6321 26638 6336 26684
rect 6382 26638 6397 26684
rect 6321 26581 6397 26638
rect 6321 26535 6336 26581
rect 6382 26535 6397 26581
rect 6321 26478 6397 26535
rect 6321 26432 6336 26478
rect 6382 26432 6397 26478
rect 6321 26375 6397 26432
rect 6321 26329 6336 26375
rect 6382 26329 6397 26375
rect 6321 26272 6397 26329
rect 6321 26226 6336 26272
rect 6382 26226 6397 26272
rect 6321 26169 6397 26226
rect 6321 26123 6336 26169
rect 6382 26123 6397 26169
rect 6321 26065 6397 26123
rect 6321 26019 6336 26065
rect 6382 26019 6397 26065
rect 6321 26006 6397 26019
rect 6565 26993 6641 27006
rect 6565 26947 6580 26993
rect 6626 26947 6641 26993
rect 6565 26890 6641 26947
rect 6565 26844 6580 26890
rect 6626 26844 6641 26890
rect 6565 26787 6641 26844
rect 6565 26741 6580 26787
rect 6626 26741 6641 26787
rect 6565 26684 6641 26741
rect 6565 26638 6580 26684
rect 6626 26638 6641 26684
rect 6565 26581 6641 26638
rect 6565 26535 6580 26581
rect 6626 26535 6641 26581
rect 6565 26478 6641 26535
rect 6565 26432 6580 26478
rect 6626 26432 6641 26478
rect 6565 26375 6641 26432
rect 6565 26329 6580 26375
rect 6626 26329 6641 26375
rect 6565 26272 6641 26329
rect 6565 26226 6580 26272
rect 6626 26226 6641 26272
rect 6565 26169 6641 26226
rect 6565 26123 6580 26169
rect 6626 26123 6641 26169
rect 6565 26065 6641 26123
rect 6565 26019 6580 26065
rect 6626 26019 6641 26065
rect 6565 25799 6641 26019
rect 6809 26993 6885 27066
rect 6809 26947 6824 26993
rect 6870 26947 6885 26993
rect 6809 26890 6885 26947
rect 6809 26844 6824 26890
rect 6870 26844 6885 26890
rect 6809 26787 6885 26844
rect 6809 26741 6824 26787
rect 6870 26741 6885 26787
rect 6809 26684 6885 26741
rect 6809 26638 6824 26684
rect 6870 26638 6885 26684
rect 6809 26581 6885 26638
rect 6809 26535 6824 26581
rect 6870 26535 6885 26581
rect 6809 26478 6885 26535
rect 6809 26432 6824 26478
rect 6870 26432 6885 26478
rect 6809 26375 6885 26432
rect 6809 26329 6824 26375
rect 6870 26329 6885 26375
rect 6809 26272 6885 26329
rect 6809 26226 6824 26272
rect 6870 26226 6885 26272
rect 6809 26169 6885 26226
rect 6809 26123 6824 26169
rect 6870 26123 6885 26169
rect 6809 26065 6885 26123
rect 6809 26019 6824 26065
rect 6870 26019 6885 26065
rect 6235 25791 6727 25799
rect 1473 25787 6759 25791
rect 1473 25735 1495 25787
rect 1651 25780 3865 25787
rect 4021 25780 6247 25787
rect 6715 25780 6759 25787
rect 1651 25735 2275 25780
rect 1473 25734 2275 25735
rect 6739 25734 6759 25780
rect 1473 25723 6759 25734
rect 6809 25617 6885 26019
rect 7053 26993 7129 27006
rect 7053 26947 7068 26993
rect 7114 26947 7129 26993
rect 7053 26890 7129 26947
rect 7053 26844 7068 26890
rect 7114 26844 7129 26890
rect 7053 26787 7129 26844
rect 7053 26741 7068 26787
rect 7114 26741 7129 26787
rect 7053 26684 7129 26741
rect 7053 26638 7068 26684
rect 7114 26638 7129 26684
rect 7053 26581 7129 26638
rect 7053 26535 7068 26581
rect 7114 26535 7129 26581
rect 7053 26478 7129 26535
rect 7053 26432 7068 26478
rect 7114 26432 7129 26478
rect 7053 26375 7129 26432
rect 7053 26329 7068 26375
rect 7114 26329 7129 26375
rect 7053 26272 7129 26329
rect 7053 26226 7068 26272
rect 7114 26226 7129 26272
rect 7053 26169 7129 26226
rect 7053 26123 7068 26169
rect 7114 26123 7129 26169
rect 7053 26065 7129 26123
rect 7053 26019 7068 26065
rect 7114 26019 7129 26065
rect 7053 25791 7129 26019
rect 7297 26993 7373 27066
rect 7297 26947 7312 26993
rect 7358 26947 7373 26993
rect 7297 26890 7373 26947
rect 7297 26844 7312 26890
rect 7358 26844 7373 26890
rect 7297 26787 7373 26844
rect 7297 26741 7312 26787
rect 7358 26741 7373 26787
rect 7297 26684 7373 26741
rect 7297 26638 7312 26684
rect 7358 26638 7373 26684
rect 7297 26581 7373 26638
rect 7297 26535 7312 26581
rect 7358 26535 7373 26581
rect 7297 26478 7373 26535
rect 7297 26432 7312 26478
rect 7358 26432 7373 26478
rect 7297 26375 7373 26432
rect 7297 26329 7312 26375
rect 7358 26329 7373 26375
rect 7297 26272 7373 26329
rect 7297 26226 7312 26272
rect 7358 26226 7373 26272
rect 7297 26169 7373 26226
rect 7297 26123 7312 26169
rect 7358 26123 7373 26169
rect 7297 26065 7373 26123
rect 7297 26019 7312 26065
rect 7358 26019 7373 26065
rect 7297 25957 7373 26019
rect 7541 26993 7617 27006
rect 7541 26947 7556 26993
rect 7602 26947 7617 26993
rect 7541 26890 7617 26947
rect 7541 26844 7556 26890
rect 7602 26844 7617 26890
rect 7541 26787 7617 26844
rect 7541 26741 7556 26787
rect 7602 26741 7617 26787
rect 7541 26684 7617 26741
rect 7541 26638 7556 26684
rect 7602 26638 7617 26684
rect 7541 26581 7617 26638
rect 7541 26535 7556 26581
rect 7602 26535 7617 26581
rect 7541 26478 7617 26535
rect 7541 26432 7556 26478
rect 7602 26432 7617 26478
rect 7541 26375 7617 26432
rect 7541 26329 7556 26375
rect 7602 26329 7617 26375
rect 7541 26272 7617 26329
rect 7541 26226 7556 26272
rect 7602 26226 7617 26272
rect 7541 26169 7617 26226
rect 7541 26123 7556 26169
rect 7602 26123 7617 26169
rect 7541 26065 7617 26123
rect 7541 26019 7556 26065
rect 7602 26019 7617 26065
rect 7541 25791 7617 26019
rect 7785 26993 7861 27066
rect 7785 26947 7800 26993
rect 7846 26947 7861 26993
rect 7785 26890 7861 26947
rect 7785 26844 7800 26890
rect 7846 26844 7861 26890
rect 7785 26787 7861 26844
rect 7785 26741 7800 26787
rect 7846 26741 7861 26787
rect 7785 26684 7861 26741
rect 7785 26638 7800 26684
rect 7846 26638 7861 26684
rect 7785 26581 7861 26638
rect 7785 26535 7800 26581
rect 7846 26535 7861 26581
rect 7785 26478 7861 26535
rect 7785 26432 7800 26478
rect 7846 26432 7861 26478
rect 7785 26375 7861 26432
rect 7785 26329 7800 26375
rect 7846 26329 7861 26375
rect 7785 26272 7861 26329
rect 7785 26226 7800 26272
rect 7846 26226 7861 26272
rect 7785 26169 7861 26226
rect 7785 26123 7800 26169
rect 7846 26123 7861 26169
rect 7785 26065 7861 26123
rect 7785 26019 7800 26065
rect 7846 26019 7861 26065
rect 7785 25957 7861 26019
rect 8029 26993 8105 27006
rect 8029 26947 8044 26993
rect 8090 26947 8105 26993
rect 8029 26890 8105 26947
rect 8029 26844 8044 26890
rect 8090 26844 8105 26890
rect 8029 26787 8105 26844
rect 8029 26741 8044 26787
rect 8090 26741 8105 26787
rect 8029 26684 8105 26741
rect 8029 26638 8044 26684
rect 8090 26638 8105 26684
rect 8029 26581 8105 26638
rect 8029 26535 8044 26581
rect 8090 26535 8105 26581
rect 8029 26478 8105 26535
rect 8029 26432 8044 26478
rect 8090 26432 8105 26478
rect 8029 26375 8105 26432
rect 8029 26329 8044 26375
rect 8090 26329 8105 26375
rect 8029 26272 8105 26329
rect 8029 26226 8044 26272
rect 8090 26226 8105 26272
rect 8029 26169 8105 26226
rect 8029 26123 8044 26169
rect 8090 26123 8105 26169
rect 8029 26065 8105 26123
rect 8029 26019 8044 26065
rect 8090 26019 8105 26065
rect 8029 25791 8105 26019
rect 10630 25888 10641 27156
rect 10687 25888 10698 27156
rect 10630 25799 10698 25888
rect 8929 25791 9109 25799
rect 10630 25791 11489 25799
rect 6935 25787 11489 25791
rect 6935 25780 8941 25787
rect 9097 25780 11311 25787
rect 6935 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25735 11311 25780
rect 11467 25735 11489 25787
rect 10687 25734 11489 25735
rect 6935 25723 11489 25734
rect 1213 25597 11749 25617
rect 1213 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11749 25597
rect 1213 25489 11749 25545
rect 1213 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11749 25489
rect 1213 25417 11749 25437
<< via1 >>
rect -309 42118 -257 45914
rect -104 45862 1092 45914
rect 1796 45862 3720 45914
rect 4166 45862 6090 45914
rect 6872 45862 8796 45914
rect 9242 45862 11166 45914
rect 11883 45862 13079 45914
rect 203 42122 1087 42174
rect 1796 42122 3720 42174
rect 4166 42122 6090 42174
rect 6872 42122 8796 42174
rect 9242 42122 11166 42174
rect 11883 42122 13079 42174
rect 13219 42118 13271 45914
rect 1495 41577 1651 41733
rect 3865 41577 4021 41733
rect 6247 41577 6715 41733
rect 8941 41577 9097 41733
rect 11311 41577 11467 41733
rect 1495 35324 1651 36000
rect 3865 35324 4021 36000
rect 6269 35946 6321 35998
rect 6393 35946 6445 35998
rect 6517 35946 6569 35998
rect 6641 35946 6693 35998
rect 6269 35822 6321 35874
rect 6393 35822 6445 35874
rect 6517 35822 6569 35874
rect 6641 35822 6693 35874
rect 6269 35698 6321 35750
rect 6393 35698 6445 35750
rect 6517 35698 6569 35750
rect 6641 35698 6693 35750
rect 6269 35574 6321 35626
rect 6393 35574 6445 35626
rect 6517 35574 6569 35626
rect 6641 35574 6693 35626
rect 6269 35450 6321 35502
rect 6393 35450 6445 35502
rect 6517 35450 6569 35502
rect 6641 35450 6693 35502
rect 6269 35326 6321 35378
rect 6393 35326 6445 35378
rect 6517 35326 6569 35378
rect 6641 35326 6693 35378
rect 8941 35324 9097 36000
rect 11311 35324 11467 36000
rect 1495 29493 1651 29649
rect 3865 29493 4021 29649
rect 6247 29493 6715 29649
rect 8941 29493 9097 29649
rect 11311 29493 11467 29649
rect 2276 29142 2328 29161
rect 2276 29034 2328 29142
rect 2276 27861 2321 29034
rect 2321 27861 2328 29034
rect 2587 28904 2639 29125
rect 2587 28858 2590 28904
rect 2590 28858 2636 28904
rect 2636 28858 2639 28904
rect 2587 28801 2639 28858
rect 2587 28755 2590 28801
rect 2590 28755 2636 28801
rect 2636 28755 2639 28801
rect 2587 28698 2639 28755
rect 2587 28652 2590 28698
rect 2590 28652 2636 28698
rect 2636 28652 2639 28698
rect 2587 28595 2639 28652
rect 2587 28549 2590 28595
rect 2590 28549 2636 28595
rect 2636 28549 2639 28595
rect 2587 28492 2639 28549
rect 2587 28446 2590 28492
rect 2590 28446 2636 28492
rect 2636 28446 2639 28492
rect 2587 28389 2639 28446
rect 2587 28343 2590 28389
rect 2590 28343 2636 28389
rect 2636 28343 2639 28389
rect 2587 28286 2639 28343
rect 2587 28240 2590 28286
rect 2590 28240 2636 28286
rect 2636 28240 2639 28286
rect 2587 28183 2639 28240
rect 2587 28137 2590 28183
rect 2590 28137 2636 28183
rect 2636 28137 2639 28183
rect 2587 28080 2639 28137
rect 2587 28034 2590 28080
rect 2590 28034 2636 28080
rect 2636 28034 2639 28080
rect 2587 27976 2639 28034
rect 2587 27930 2590 27976
rect 2590 27930 2636 27976
rect 2636 27930 2639 27976
rect 2587 27929 2639 27930
rect 3075 28904 3127 29125
rect 3075 28858 3078 28904
rect 3078 28858 3124 28904
rect 3124 28858 3127 28904
rect 3075 28801 3127 28858
rect 3075 28755 3078 28801
rect 3078 28755 3124 28801
rect 3124 28755 3127 28801
rect 3075 28698 3127 28755
rect 3075 28652 3078 28698
rect 3078 28652 3124 28698
rect 3124 28652 3127 28698
rect 3075 28595 3127 28652
rect 3075 28549 3078 28595
rect 3078 28549 3124 28595
rect 3124 28549 3127 28595
rect 3075 28492 3127 28549
rect 3075 28446 3078 28492
rect 3078 28446 3124 28492
rect 3124 28446 3127 28492
rect 3075 28389 3127 28446
rect 3075 28343 3078 28389
rect 3078 28343 3124 28389
rect 3124 28343 3127 28389
rect 3075 28286 3127 28343
rect 3075 28240 3078 28286
rect 3078 28240 3124 28286
rect 3124 28240 3127 28286
rect 3075 28183 3127 28240
rect 3075 28137 3078 28183
rect 3078 28137 3124 28183
rect 3124 28137 3127 28183
rect 3075 28080 3127 28137
rect 3075 28034 3078 28080
rect 3078 28034 3124 28080
rect 3124 28034 3127 28080
rect 3075 27976 3127 28034
rect 3075 27930 3078 27976
rect 3078 27930 3124 27976
rect 3124 27930 3127 27976
rect 3075 27929 3127 27930
rect 3563 28904 3615 29125
rect 3563 28858 3566 28904
rect 3566 28858 3612 28904
rect 3612 28858 3615 28904
rect 3563 28801 3615 28858
rect 3563 28755 3566 28801
rect 3566 28755 3612 28801
rect 3612 28755 3615 28801
rect 3563 28698 3615 28755
rect 3563 28652 3566 28698
rect 3566 28652 3612 28698
rect 3612 28652 3615 28698
rect 3563 28595 3615 28652
rect 3563 28549 3566 28595
rect 3566 28549 3612 28595
rect 3612 28549 3615 28595
rect 3563 28492 3615 28549
rect 3563 28446 3566 28492
rect 3566 28446 3612 28492
rect 3612 28446 3615 28492
rect 3563 28389 3615 28446
rect 3563 28343 3566 28389
rect 3566 28343 3612 28389
rect 3612 28343 3615 28389
rect 3563 28286 3615 28343
rect 3563 28240 3566 28286
rect 3566 28240 3612 28286
rect 3612 28240 3615 28286
rect 3563 28183 3615 28240
rect 3563 28137 3566 28183
rect 3566 28137 3612 28183
rect 3612 28137 3615 28183
rect 3563 28080 3615 28137
rect 3563 28034 3566 28080
rect 3566 28034 3612 28080
rect 3612 28034 3615 28080
rect 3563 27976 3615 28034
rect 3563 27930 3566 27976
rect 3566 27930 3612 27976
rect 3612 27930 3615 27976
rect 3563 27929 3615 27930
rect 4467 28904 4519 29125
rect 4467 28858 4470 28904
rect 4470 28858 4516 28904
rect 4516 28858 4519 28904
rect 4467 28801 4519 28858
rect 4467 28755 4470 28801
rect 4470 28755 4516 28801
rect 4516 28755 4519 28801
rect 4467 28698 4519 28755
rect 4467 28652 4470 28698
rect 4470 28652 4516 28698
rect 4516 28652 4519 28698
rect 4467 28595 4519 28652
rect 4467 28549 4470 28595
rect 4470 28549 4516 28595
rect 4516 28549 4519 28595
rect 4467 28492 4519 28549
rect 4467 28446 4470 28492
rect 4470 28446 4516 28492
rect 4516 28446 4519 28492
rect 4467 28389 4519 28446
rect 4467 28343 4470 28389
rect 4470 28343 4516 28389
rect 4516 28343 4519 28389
rect 4467 28286 4519 28343
rect 4467 28240 4470 28286
rect 4470 28240 4516 28286
rect 4516 28240 4519 28286
rect 4467 28183 4519 28240
rect 4467 28137 4470 28183
rect 4470 28137 4516 28183
rect 4516 28137 4519 28183
rect 4467 28080 4519 28137
rect 4467 28034 4470 28080
rect 4470 28034 4516 28080
rect 4516 28034 4519 28080
rect 4467 27976 4519 28034
rect 4467 27930 4470 27976
rect 4470 27930 4516 27976
rect 4516 27930 4519 27976
rect 4467 27929 4519 27930
rect 4955 28904 5007 29125
rect 4955 28858 4958 28904
rect 4958 28858 5004 28904
rect 5004 28858 5007 28904
rect 4955 28801 5007 28858
rect 4955 28755 4958 28801
rect 4958 28755 5004 28801
rect 5004 28755 5007 28801
rect 4955 28698 5007 28755
rect 4955 28652 4958 28698
rect 4958 28652 5004 28698
rect 5004 28652 5007 28698
rect 4955 28595 5007 28652
rect 4955 28549 4958 28595
rect 4958 28549 5004 28595
rect 5004 28549 5007 28595
rect 4955 28492 5007 28549
rect 4955 28446 4958 28492
rect 4958 28446 5004 28492
rect 5004 28446 5007 28492
rect 4955 28389 5007 28446
rect 4955 28343 4958 28389
rect 4958 28343 5004 28389
rect 5004 28343 5007 28389
rect 4955 28286 5007 28343
rect 4955 28240 4958 28286
rect 4958 28240 5004 28286
rect 5004 28240 5007 28286
rect 4955 28183 5007 28240
rect 4955 28137 4958 28183
rect 4958 28137 5004 28183
rect 5004 28137 5007 28183
rect 4955 28080 5007 28137
rect 4955 28034 4958 28080
rect 4958 28034 5004 28080
rect 5004 28034 5007 28080
rect 4955 27976 5007 28034
rect 4955 27930 4958 27976
rect 4958 27930 5004 27976
rect 5004 27930 5007 27976
rect 4955 27929 5007 27930
rect 5443 28904 5495 29125
rect 5443 28858 5446 28904
rect 5446 28858 5492 28904
rect 5492 28858 5495 28904
rect 5443 28801 5495 28858
rect 5443 28755 5446 28801
rect 5446 28755 5492 28801
rect 5492 28755 5495 28801
rect 5443 28698 5495 28755
rect 5443 28652 5446 28698
rect 5446 28652 5492 28698
rect 5492 28652 5495 28698
rect 5443 28595 5495 28652
rect 5443 28549 5446 28595
rect 5446 28549 5492 28595
rect 5492 28549 5495 28595
rect 5443 28492 5495 28549
rect 5443 28446 5446 28492
rect 5446 28446 5492 28492
rect 5492 28446 5495 28492
rect 5443 28389 5495 28446
rect 5443 28343 5446 28389
rect 5446 28343 5492 28389
rect 5492 28343 5495 28389
rect 5443 28286 5495 28343
rect 5443 28240 5446 28286
rect 5446 28240 5492 28286
rect 5492 28240 5495 28286
rect 5443 28183 5495 28240
rect 5443 28137 5446 28183
rect 5446 28137 5492 28183
rect 5492 28137 5495 28183
rect 5443 28080 5495 28137
rect 5443 28034 5446 28080
rect 5446 28034 5492 28080
rect 5492 28034 5495 28080
rect 5443 27976 5495 28034
rect 5443 27930 5446 27976
rect 5446 27930 5492 27976
rect 5492 27930 5495 27976
rect 5443 27929 5495 27930
rect 5931 28904 5983 29125
rect 5931 28858 5934 28904
rect 5934 28858 5980 28904
rect 5980 28858 5983 28904
rect 5931 28801 5983 28858
rect 5931 28755 5934 28801
rect 5934 28755 5980 28801
rect 5980 28755 5983 28801
rect 5931 28698 5983 28755
rect 5931 28652 5934 28698
rect 5934 28652 5980 28698
rect 5980 28652 5983 28698
rect 5931 28595 5983 28652
rect 5931 28549 5934 28595
rect 5934 28549 5980 28595
rect 5980 28549 5983 28595
rect 5931 28492 5983 28549
rect 5931 28446 5934 28492
rect 5934 28446 5980 28492
rect 5980 28446 5983 28492
rect 5931 28389 5983 28446
rect 5931 28343 5934 28389
rect 5934 28343 5980 28389
rect 5980 28343 5983 28389
rect 5931 28286 5983 28343
rect 5931 28240 5934 28286
rect 5934 28240 5980 28286
rect 5980 28240 5983 28286
rect 5931 28183 5983 28240
rect 5931 28137 5934 28183
rect 5934 28137 5980 28183
rect 5980 28137 5983 28183
rect 5931 28080 5983 28137
rect 5931 28034 5934 28080
rect 5934 28034 5980 28080
rect 5980 28034 5983 28080
rect 5931 27976 5983 28034
rect 5931 27930 5934 27976
rect 5934 27930 5980 27976
rect 5980 27930 5983 27976
rect 5931 27929 5983 27930
rect 6907 28904 6959 29125
rect 6907 28858 6910 28904
rect 6910 28858 6956 28904
rect 6956 28858 6959 28904
rect 6907 28801 6959 28858
rect 6907 28755 6910 28801
rect 6910 28755 6956 28801
rect 6956 28755 6959 28801
rect 6907 28698 6959 28755
rect 6907 28652 6910 28698
rect 6910 28652 6956 28698
rect 6956 28652 6959 28698
rect 6907 28595 6959 28652
rect 6907 28549 6910 28595
rect 6910 28549 6956 28595
rect 6956 28549 6959 28595
rect 6907 28492 6959 28549
rect 6907 28446 6910 28492
rect 6910 28446 6956 28492
rect 6956 28446 6959 28492
rect 6907 28389 6959 28446
rect 6907 28343 6910 28389
rect 6910 28343 6956 28389
rect 6956 28343 6959 28389
rect 6907 28286 6959 28343
rect 6907 28240 6910 28286
rect 6910 28240 6956 28286
rect 6956 28240 6959 28286
rect 6907 28183 6959 28240
rect 6907 28137 6910 28183
rect 6910 28137 6956 28183
rect 6956 28137 6959 28183
rect 6907 28080 6959 28137
rect 6907 28034 6910 28080
rect 6910 28034 6956 28080
rect 6956 28034 6959 28080
rect 6907 27976 6959 28034
rect 6907 27930 6910 27976
rect 6910 27930 6956 27976
rect 6956 27930 6959 27976
rect 6907 27929 6959 27930
rect 7395 28904 7447 29125
rect 7395 28858 7398 28904
rect 7398 28858 7444 28904
rect 7444 28858 7447 28904
rect 7395 28801 7447 28858
rect 7395 28755 7398 28801
rect 7398 28755 7444 28801
rect 7444 28755 7447 28801
rect 7395 28698 7447 28755
rect 7395 28652 7398 28698
rect 7398 28652 7444 28698
rect 7444 28652 7447 28698
rect 7395 28595 7447 28652
rect 7395 28549 7398 28595
rect 7398 28549 7444 28595
rect 7444 28549 7447 28595
rect 7395 28492 7447 28549
rect 7395 28446 7398 28492
rect 7398 28446 7444 28492
rect 7444 28446 7447 28492
rect 7395 28389 7447 28446
rect 7395 28343 7398 28389
rect 7398 28343 7444 28389
rect 7444 28343 7447 28389
rect 7395 28286 7447 28343
rect 7395 28240 7398 28286
rect 7398 28240 7444 28286
rect 7444 28240 7447 28286
rect 7395 28183 7447 28240
rect 7395 28137 7398 28183
rect 7398 28137 7444 28183
rect 7444 28137 7447 28183
rect 7395 28080 7447 28137
rect 7395 28034 7398 28080
rect 7398 28034 7444 28080
rect 7444 28034 7447 28080
rect 7395 27976 7447 28034
rect 7395 27930 7398 27976
rect 7398 27930 7444 27976
rect 7444 27930 7447 27976
rect 7395 27929 7447 27930
rect 7883 28904 7935 29125
rect 7883 28858 7886 28904
rect 7886 28858 7932 28904
rect 7932 28858 7935 28904
rect 7883 28801 7935 28858
rect 7883 28755 7886 28801
rect 7886 28755 7932 28801
rect 7932 28755 7935 28801
rect 7883 28698 7935 28755
rect 7883 28652 7886 28698
rect 7886 28652 7932 28698
rect 7932 28652 7935 28698
rect 7883 28595 7935 28652
rect 7883 28549 7886 28595
rect 7886 28549 7932 28595
rect 7932 28549 7935 28595
rect 7883 28492 7935 28549
rect 7883 28446 7886 28492
rect 7886 28446 7932 28492
rect 7932 28446 7935 28492
rect 7883 28389 7935 28446
rect 7883 28343 7886 28389
rect 7886 28343 7932 28389
rect 7932 28343 7935 28389
rect 7883 28286 7935 28343
rect 7883 28240 7886 28286
rect 7886 28240 7932 28286
rect 7932 28240 7935 28286
rect 7883 28183 7935 28240
rect 7883 28137 7886 28183
rect 7886 28137 7932 28183
rect 7932 28137 7935 28183
rect 7883 28080 7935 28137
rect 7883 28034 7886 28080
rect 7886 28034 7932 28080
rect 7932 28034 7935 28080
rect 7883 27976 7935 28034
rect 7883 27930 7886 27976
rect 7886 27930 7932 27976
rect 7932 27930 7935 27976
rect 7883 27929 7935 27930
rect 8371 28904 8423 29125
rect 8371 28858 8374 28904
rect 8374 28858 8420 28904
rect 8420 28858 8423 28904
rect 8371 28801 8423 28858
rect 8371 28755 8374 28801
rect 8374 28755 8420 28801
rect 8420 28755 8423 28801
rect 8371 28698 8423 28755
rect 8371 28652 8374 28698
rect 8374 28652 8420 28698
rect 8420 28652 8423 28698
rect 8371 28595 8423 28652
rect 8371 28549 8374 28595
rect 8374 28549 8420 28595
rect 8420 28549 8423 28595
rect 8371 28492 8423 28549
rect 8371 28446 8374 28492
rect 8374 28446 8420 28492
rect 8420 28446 8423 28492
rect 8371 28389 8423 28446
rect 8371 28343 8374 28389
rect 8374 28343 8420 28389
rect 8420 28343 8423 28389
rect 8371 28286 8423 28343
rect 8371 28240 8374 28286
rect 8374 28240 8420 28286
rect 8420 28240 8423 28286
rect 8371 28183 8423 28240
rect 8371 28137 8374 28183
rect 8374 28137 8420 28183
rect 8420 28137 8423 28183
rect 8371 28080 8423 28137
rect 8371 28034 8374 28080
rect 8374 28034 8420 28080
rect 8420 28034 8423 28080
rect 8371 27976 8423 28034
rect 8371 27930 8374 27976
rect 8374 27930 8420 27976
rect 8420 27930 8423 27976
rect 8371 27929 8423 27930
rect 9347 28904 9399 29125
rect 9347 28858 9350 28904
rect 9350 28858 9396 28904
rect 9396 28858 9399 28904
rect 9347 28801 9399 28858
rect 9347 28755 9350 28801
rect 9350 28755 9396 28801
rect 9396 28755 9399 28801
rect 9347 28698 9399 28755
rect 9347 28652 9350 28698
rect 9350 28652 9396 28698
rect 9396 28652 9399 28698
rect 9347 28595 9399 28652
rect 9347 28549 9350 28595
rect 9350 28549 9396 28595
rect 9396 28549 9399 28595
rect 9347 28492 9399 28549
rect 9347 28446 9350 28492
rect 9350 28446 9396 28492
rect 9396 28446 9399 28492
rect 9347 28389 9399 28446
rect 9347 28343 9350 28389
rect 9350 28343 9396 28389
rect 9396 28343 9399 28389
rect 9347 28286 9399 28343
rect 9347 28240 9350 28286
rect 9350 28240 9396 28286
rect 9396 28240 9399 28286
rect 9347 28183 9399 28240
rect 9347 28137 9350 28183
rect 9350 28137 9396 28183
rect 9396 28137 9399 28183
rect 9347 28080 9399 28137
rect 9347 28034 9350 28080
rect 9350 28034 9396 28080
rect 9396 28034 9399 28080
rect 9347 27976 9399 28034
rect 9347 27930 9350 27976
rect 9350 27930 9396 27976
rect 9396 27930 9399 27976
rect 9347 27929 9399 27930
rect 9835 28904 9887 29125
rect 9835 28858 9838 28904
rect 9838 28858 9884 28904
rect 9884 28858 9887 28904
rect 9835 28801 9887 28858
rect 9835 28755 9838 28801
rect 9838 28755 9884 28801
rect 9884 28755 9887 28801
rect 9835 28698 9887 28755
rect 9835 28652 9838 28698
rect 9838 28652 9884 28698
rect 9884 28652 9887 28698
rect 9835 28595 9887 28652
rect 9835 28549 9838 28595
rect 9838 28549 9884 28595
rect 9884 28549 9887 28595
rect 9835 28492 9887 28549
rect 9835 28446 9838 28492
rect 9838 28446 9884 28492
rect 9884 28446 9887 28492
rect 9835 28389 9887 28446
rect 9835 28343 9838 28389
rect 9838 28343 9884 28389
rect 9884 28343 9887 28389
rect 9835 28286 9887 28343
rect 9835 28240 9838 28286
rect 9838 28240 9884 28286
rect 9884 28240 9887 28286
rect 9835 28183 9887 28240
rect 9835 28137 9838 28183
rect 9838 28137 9884 28183
rect 9884 28137 9887 28183
rect 9835 28080 9887 28137
rect 9835 28034 9838 28080
rect 9838 28034 9884 28080
rect 9884 28034 9887 28080
rect 9835 27976 9887 28034
rect 9835 27930 9838 27976
rect 9838 27930 9884 27976
rect 9884 27930 9887 27976
rect 9835 27929 9887 27930
rect 10323 28904 10375 29125
rect 10323 28858 10326 28904
rect 10326 28858 10372 28904
rect 10372 28858 10375 28904
rect 10323 28801 10375 28858
rect 10323 28755 10326 28801
rect 10326 28755 10372 28801
rect 10372 28755 10375 28801
rect 10323 28698 10375 28755
rect 10323 28652 10326 28698
rect 10326 28652 10372 28698
rect 10372 28652 10375 28698
rect 10323 28595 10375 28652
rect 10323 28549 10326 28595
rect 10326 28549 10372 28595
rect 10372 28549 10375 28595
rect 10323 28492 10375 28549
rect 10323 28446 10326 28492
rect 10326 28446 10372 28492
rect 10372 28446 10375 28492
rect 10323 28389 10375 28446
rect 10323 28343 10326 28389
rect 10326 28343 10372 28389
rect 10372 28343 10375 28389
rect 10323 28286 10375 28343
rect 10323 28240 10326 28286
rect 10326 28240 10372 28286
rect 10372 28240 10375 28286
rect 10323 28183 10375 28240
rect 10323 28137 10326 28183
rect 10326 28137 10372 28183
rect 10372 28137 10375 28183
rect 10323 28080 10375 28137
rect 10323 28034 10326 28080
rect 10326 28034 10372 28080
rect 10372 28034 10375 28080
rect 10323 27976 10375 28034
rect 10323 27930 10326 27976
rect 10326 27930 10372 27976
rect 10372 27930 10375 27976
rect 10323 27929 10375 27930
rect 10634 29034 10686 29125
rect 10634 27929 10641 29034
rect 10641 27929 10686 29034
rect 3865 27439 4021 27484
rect 6257 27439 6517 27484
rect 3865 27432 4021 27439
rect 6257 27432 6517 27439
rect 8941 27439 9097 27484
rect 8941 27432 9097 27439
rect 1495 25735 1651 25787
rect 3865 25780 4021 25787
rect 6247 25780 6715 25787
rect 3865 25735 4021 25780
rect 6247 25735 6715 25780
rect 8941 25780 9097 25787
rect 8941 25735 9097 25780
rect 11311 25735 11467 25787
rect 1233 25545 1285 25597
rect 1341 25545 1393 25597
rect 11569 25545 11621 25597
rect 11677 25545 11729 25597
rect 1233 25437 1285 25489
rect 1341 25437 1393 25489
rect 11569 25437 11621 25489
rect 11677 25437 11729 25489
<< metal2 >>
rect -747 45914 1153 46134
rect -747 42118 -309 45914
rect -257 45862 -104 45914
rect 1092 45862 1153 45914
rect -257 42174 1153 45862
rect -257 42122 203 42174
rect 1087 42122 1153 42174
rect -257 42118 1153 42122
rect -747 25617 1153 42118
rect 1473 41733 1673 46134
rect 1473 41577 1495 41733
rect 1651 41577 1673 41733
rect 1473 36000 1673 41577
rect 1473 35324 1495 36000
rect 1651 35324 1673 36000
rect 1473 29649 1673 35324
rect 1473 29493 1495 29649
rect 1651 29493 1673 29649
rect 1473 25787 1673 29493
rect 1473 25735 1495 25787
rect 1651 25735 1673 25787
rect 1473 25617 1673 25735
rect 1733 45914 3783 46134
rect 1733 45862 1796 45914
rect 3720 45862 3783 45914
rect 1733 42174 3783 45862
rect 1733 42122 1796 42174
rect 3720 42122 3783 42174
rect 1733 29161 3783 42122
rect 1733 27861 2276 29161
rect 2328 29125 3783 29161
rect 2328 27929 2587 29125
rect 2639 27929 3075 29125
rect 3127 27929 3563 29125
rect 3615 27929 3783 29125
rect 2328 27861 3783 27929
rect 1733 25617 3783 27861
rect 3843 41733 4043 46134
rect 3843 41577 3865 41733
rect 4021 41577 4043 41733
rect 3843 36000 4043 41577
rect 3843 35324 3865 36000
rect 4021 35324 4043 36000
rect 3843 29649 4043 35324
rect 3843 29493 3865 29649
rect 4021 29493 4043 29649
rect 3843 27484 4043 29493
rect 3843 27432 3865 27484
rect 4021 27432 4043 27484
rect 3843 25787 4043 27432
rect 3843 25735 3865 25787
rect 4021 25735 4043 25787
rect 3843 25617 4043 25735
rect 4103 45914 6153 46134
rect 4103 45862 4166 45914
rect 6090 45862 6153 45914
rect 4103 42174 6153 45862
rect 4103 42122 4166 42174
rect 6090 42122 6153 42174
rect 4103 29125 6153 42122
rect 4103 27929 4467 29125
rect 4519 27929 4955 29125
rect 5007 27929 5443 29125
rect 5495 27929 5931 29125
rect 5983 27929 6153 29125
rect 4103 25617 6153 27929
rect 6213 41733 6749 46134
rect 6213 41577 6247 41733
rect 6715 41577 6749 41733
rect 6213 35998 6749 41577
rect 6213 35946 6269 35998
rect 6321 35946 6393 35998
rect 6445 35946 6517 35998
rect 6569 35946 6641 35998
rect 6693 35946 6749 35998
rect 6213 35874 6749 35946
rect 6213 35822 6269 35874
rect 6321 35822 6393 35874
rect 6445 35822 6517 35874
rect 6569 35822 6641 35874
rect 6693 35822 6749 35874
rect 6213 35750 6749 35822
rect 6213 35698 6269 35750
rect 6321 35698 6393 35750
rect 6445 35698 6517 35750
rect 6569 35698 6641 35750
rect 6693 35698 6749 35750
rect 6213 35626 6749 35698
rect 6213 35574 6269 35626
rect 6321 35574 6393 35626
rect 6445 35574 6517 35626
rect 6569 35574 6641 35626
rect 6693 35574 6749 35626
rect 6213 35502 6749 35574
rect 6213 35450 6269 35502
rect 6321 35450 6393 35502
rect 6445 35450 6517 35502
rect 6569 35450 6641 35502
rect 6693 35450 6749 35502
rect 6213 35378 6749 35450
rect 6213 35326 6269 35378
rect 6321 35326 6393 35378
rect 6445 35326 6517 35378
rect 6569 35326 6641 35378
rect 6693 35326 6749 35378
rect 6213 29649 6749 35326
rect 6213 29493 6247 29649
rect 6715 29493 6749 29649
rect 6213 27484 6749 29493
rect 6213 27432 6257 27484
rect 6517 27432 6749 27484
rect 6213 25787 6749 27432
rect 6213 25735 6247 25787
rect 6715 25735 6749 25787
rect 6213 25617 6749 25735
rect 6809 45914 8859 46134
rect 6809 45862 6872 45914
rect 8796 45862 8859 45914
rect 6809 42174 8859 45862
rect 6809 42122 6872 42174
rect 8796 42122 8859 42174
rect 6809 29125 8859 42122
rect 6809 27929 6907 29125
rect 6959 27929 7395 29125
rect 7447 27929 7883 29125
rect 7935 27929 8371 29125
rect 8423 27929 8859 29125
rect 6809 25617 8859 27929
rect 8919 41733 9119 46134
rect 8919 41577 8941 41733
rect 9097 41577 9119 41733
rect 8919 36000 9119 41577
rect 8919 35324 8941 36000
rect 9097 35324 9119 36000
rect 8919 29649 9119 35324
rect 8919 29493 8941 29649
rect 9097 29493 9119 29649
rect 8919 27484 9119 29493
rect 8919 27432 8941 27484
rect 9097 27432 9119 27484
rect 8919 25787 9119 27432
rect 8919 25735 8941 25787
rect 9097 25735 9119 25787
rect 8919 25617 9119 25735
rect 9179 45914 11229 46134
rect 9179 45862 9242 45914
rect 11166 45862 11229 45914
rect 9179 42174 11229 45862
rect 9179 42122 9242 42174
rect 11166 42122 11229 42174
rect 9179 29125 11229 42122
rect 9179 27929 9347 29125
rect 9399 27929 9835 29125
rect 9887 27929 10323 29125
rect 10375 27929 10634 29125
rect 10686 27929 11229 29125
rect 9179 25617 11229 27929
rect 11289 41733 11489 46134
rect 11289 41577 11311 41733
rect 11467 41577 11489 41733
rect 11289 36000 11489 41577
rect 11289 35324 11311 36000
rect 11467 35324 11489 36000
rect 11289 29649 11489 35324
rect 11289 29493 11311 29649
rect 11467 29493 11489 29649
rect 11289 25787 11489 29493
rect 11289 25735 11311 25787
rect 11467 25735 11489 25787
rect 11289 25617 11489 25735
rect 11809 45914 13709 46134
rect 11809 45862 11883 45914
rect 13079 45862 13219 45914
rect 11809 42174 13219 45862
rect 11809 42122 11883 42174
rect 13079 42122 13219 42174
rect 11809 42118 13219 42122
rect 13271 42118 13709 45914
rect 11809 25617 13709 42118
rect 1221 25597 1405 25609
rect 1221 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 1405 25597
rect 1221 25489 1405 25545
rect 1221 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 1405 25489
rect 1221 25425 1405 25437
rect 11557 25597 11741 25609
rect 11557 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11741 25597
rect 11557 25489 11741 25545
rect 11557 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11741 25489
rect 11557 25425 11741 25437
use M1_NWELL_CDNS_40661953145107  M1_NWELL_CDNS_40661953145107_0
timestamp 1666464484
transform 1 0 6481 0 1 29165
box 0 0 1 1
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_0
timestamp 1666464484
transform 1 0 10664 0 1 28447
box 0 0 1 1
use M1_NWELL_CDNS_40661953145111  M1_NWELL_CDNS_40661953145111_1
timestamp 1666464484
transform 1 0 2298 0 1 28447
box 0 0 1 1
use M1_POLY2_CDNS_40661953145105  M1_POLY2_CDNS_40661953145105_0
timestamp 1666464484
transform 1 0 3101 0 1 27687
box 0 0 1 1
use M1_POLY2_CDNS_40661953145106  M1_POLY2_CDNS_40661953145106_0
timestamp 1666464484
transform 1 0 4142 0 1 27108
box 0 0 1 1
use M1_POLY2_CDNS_40661953145108  M1_POLY2_CDNS_40661953145108_0
timestamp 1666464484
transform 1 0 3955 0 1 27687
box 0 0 1 1
use M1_POLY2_CDNS_40661953145109  M1_POLY2_CDNS_40661953145109_0
timestamp 1666464484
transform 1 0 7335 0 1 27236
box 0 0 1 1
use M1_POLY2_CDNS_40661953145109  M1_POLY2_CDNS_40661953145109_1
timestamp 1666464484
transform 1 0 5871 0 1 27236
box 0 0 1 1
use M1_POLY2_CDNS_40661953145110  M1_POLY2_CDNS_40661953145110_0
timestamp 1666464484
transform 1 0 7421 0 1 27687
box 0 0 1 1
use M1_PSUB_CDNS_40661953145102  M1_PSUB_CDNS_40661953145102_0
timestamp 1666464484
transform 1 0 10664 0 -1 26522
box 0 0 1 1
use M1_PSUB_CDNS_40661953145102  M1_PSUB_CDNS_40661953145102_1
timestamp 1666464484
transform 1 0 2298 0 -1 26522
box 0 0 1 1
use M1_PSUB_CDNS_40661953145123  M1_PSUB_CDNS_40661953145123_0
timestamp 1666464484
transform 1 0 5132 0 1 27462
box 0 0 1 1
use M1_PSUB_CDNS_40661953145124  M1_PSUB_CDNS_40661953145124_0
timestamp 1666464484
transform 1 0 8555 0 1 27462
box 0 0 1 1
use M2_M1_CDNS_40661953145103  M2_M1_CDNS_40661953145103_0
timestamp 1666464484
transform 1 0 11649 0 1 25517
box 0 0 1 1
use M2_M1_CDNS_40661953145103  M2_M1_CDNS_40661953145103_1
timestamp 1666464484
transform 1 0 1313 0 1 25517
box 0 0 1 1
use M2_M1_CDNS_40661953145104  M2_M1_CDNS_40661953145104_0
timestamp 1666464484
transform 1 0 6481 0 1 41655
box 0 0 1 1
use M2_M1_CDNS_40661953145104  M2_M1_CDNS_40661953145104_1
timestamp 1666464484
transform 1 0 6481 0 1 29571
box 0 0 1 1
use M2_M1_CDNS_40661953145112  M2_M1_CDNS_40661953145112_0
timestamp 1666464484
transform -1 0 6481 0 1 25761
box 0 0 1 1
use M2_M1_CDNS_40661953145113  M2_M1_CDNS_40661953145113_0
timestamp 1666464484
transform 1 0 645 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145114  M2_M1_CDNS_40661953145114_0
timestamp 1666464484
transform 1 0 12481 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145114  M2_M1_CDNS_40661953145114_1
timestamp 1666464484
transform 1 0 12481 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145114  M2_M1_CDNS_40661953145114_2
timestamp 1666464484
transform 1 0 494 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_0
timestamp 1666464484
transform 1 0 1573 0 1 41655
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_1
timestamp 1666464484
transform 1 0 1573 0 1 29571
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_2
timestamp 1666464484
transform 1 0 3943 0 1 29571
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_3
timestamp 1666464484
transform 1 0 11389 0 1 29571
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_4
timestamp 1666464484
transform 1 0 3943 0 1 41655
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_5
timestamp 1666464484
transform 1 0 9019 0 1 29571
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_6
timestamp 1666464484
transform 1 0 9019 0 1 41655
box 0 0 1 1
use M2_M1_CDNS_40661953145115  M2_M1_CDNS_40661953145115_7
timestamp 1666464484
transform 1 0 11389 0 1 41655
box 0 0 1 1
use M2_M1_CDNS_40661953145116  M2_M1_CDNS_40661953145116_0
timestamp 1666464484
transform 1 0 13245 0 1 44016
box 0 0 1 1
use M2_M1_CDNS_40661953145116  M2_M1_CDNS_40661953145116_1
timestamp 1666464484
transform 1 0 -283 0 1 44016
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_0
timestamp 1666464484
transform -1 0 3943 0 1 25761
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_1
timestamp 1666464484
transform -1 0 11389 0 1 25761
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_2
timestamp 1666464484
transform -1 0 9019 0 1 25761
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_3
timestamp 1666464484
transform -1 0 9019 0 1 27458
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_4
timestamp 1666464484
transform -1 0 3943 0 1 27458
box 0 0 1 1
use M2_M1_CDNS_40661953145117  M2_M1_CDNS_40661953145117_5
timestamp 1666464484
transform 1 0 1573 0 1 25761
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_0
timestamp 1666464484
transform 1 0 2758 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_1
timestamp 1666464484
transform 1 0 2758 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_2
timestamp 1666464484
transform 1 0 5128 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_3
timestamp 1666464484
transform 1 0 5128 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_4
timestamp 1666464484
transform 1 0 7834 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_5
timestamp 1666464484
transform 1 0 7834 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_6
timestamp 1666464484
transform 1 0 10204 0 1 42148
box 0 0 1 1
use M2_M1_CDNS_40661953145118  M2_M1_CDNS_40661953145118_7
timestamp 1666464484
transform 1 0 10204 0 1 45888
box 0 0 1 1
use M2_M1_CDNS_40661953145119  M2_M1_CDNS_40661953145119_0
timestamp 1666464484
transform 1 0 11389 0 1 35662
box 0 0 1 1
use M2_M1_CDNS_40661953145119  M2_M1_CDNS_40661953145119_1
timestamp 1666464484
transform 1 0 9019 0 1 35662
box 0 0 1 1
use M2_M1_CDNS_40661953145119  M2_M1_CDNS_40661953145119_2
timestamp 1666464484
transform 1 0 3943 0 1 35662
box 0 0 1 1
use M2_M1_CDNS_40661953145119  M2_M1_CDNS_40661953145119_3
timestamp 1666464484
transform 1 0 1573 0 1 35662
box 0 0 1 1
use M2_M1_CDNS_40661953145120  M2_M1_CDNS_40661953145120_0
timestamp 1666464484
transform 1 0 2302 0 1 28511
box 0 0 1 1
use M2_M1_CDNS_40661953145121  M2_M1_CDNS_40661953145121_0
timestamp 1666464484
transform 1 0 6481 0 1 35662
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_0
timestamp 1666464484
transform 1 0 5957 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_1
timestamp 1666464484
transform 1 0 5469 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_2
timestamp 1666464484
transform 1 0 4981 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_3
timestamp 1666464484
transform 1 0 4493 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_4
timestamp 1666464484
transform 1 0 3589 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_5
timestamp 1666464484
transform 1 0 3101 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_6
timestamp 1666464484
transform 1 0 2613 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_7
timestamp 1666464484
transform 1 0 6933 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_8
timestamp 1666464484
transform 1 0 7909 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_9
timestamp 1666464484
transform 1 0 8397 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_10
timestamp 1666464484
transform 1 0 9373 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_11
timestamp 1666464484
transform 1 0 9861 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_12
timestamp 1666464484
transform 1 0 10349 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_13
timestamp 1666464484
transform 1 0 10660 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145122  M2_M1_CDNS_40661953145122_14
timestamp 1666464484
transform 1 0 7421 0 1 28527
box 0 0 1 1
use M2_M1_CDNS_40661953145125  M2_M1_CDNS_40661953145125_0
timestamp 1666464484
transform -1 0 6387 0 1 27458
box 0 0 1 1
use comp018green_esd_rc_v5p0  comp018green_esd_rc_v5p0_0
timestamp 1666464484
transform 1 0 -356 0 -1 46507
box -51 491 13725 17038
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_0
timestamp 1666464484
transform 1 0 6655 0 1 26006
box 0 0 1 1
use nmos_6p0_CDNS_406619531458  nmos_6p0_CDNS_406619531458_1
timestamp 1666464484
transform 1 0 5191 0 1 26006
box 0 0 1 1
use nmos_6p0_CDNS_406619531459  nmos_6p0_CDNS_406619531459_0
timestamp 1666464484
transform 1 0 4129 0 1 26006
box 0 0 1 1
use nmos_clamp_20_50_4_DVDD  nmos_clamp_20_50_4_DVDD_0
timestamp 1666464484
transform 1 0 0 0 1 0
box -747 -51 13709 25617
use pmos_6p0_CDNS_406619531452  pmos_6p0_CDNS_406619531452_0
timestamp 1666464484
transform 1 0 2665 0 1 27917
box 0 0 1 1
use pmos_6p0_CDNS_406619531455  pmos_6p0_CDNS_406619531455_0
timestamp 1666464484
transform 1 0 4545 0 1 27917
box 0 0 1 1
use pmos_6p0_CDNS_406619531456  pmos_6p0_CDNS_406619531456_0
timestamp 1666464484
transform 1 0 3641 0 1 27917
box 0 0 1 1
<< properties >>
string GDS_END 2009734
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 1992714
string path 287.225 644.025 265.750 644.025 
<< end >>
