magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 227 88 300
rect 193 227 312 300
rect 417 227 536 300
rect 641 227 760 300
rect 865 227 984 300
rect -31 -74 88 -1
rect 193 -74 312 -1
rect 417 -74 536 -1
rect 641 -74 760 -1
rect 865 -74 984 -1
use nmos_5p04310590878134_256x8m81  nmos_5p04310590878134_256x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 1104 272
<< properties >>
string GDS_END 351898
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 351136
<< end >>
