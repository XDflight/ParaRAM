magic
tech gf180mcuB
timestamp 1666464484
<< metal1 >>
rect 0 147 62 159
rect 11 106 16 147
rect 28 86 33 140
rect 45 106 50 147
rect 26 80 36 86
rect 12 67 22 73
rect 28 40 33 80
rect 38 54 48 60
rect 14 35 33 40
rect 14 16 19 35
rect 42 9 47 33
rect 0 -3 62 9
<< metal2 >>
rect 10 154 18 155
rect 34 154 42 155
rect 9 148 19 154
rect 33 148 43 154
rect 10 147 18 148
rect 34 147 42 148
rect 26 79 36 87
rect 12 66 22 74
rect 38 53 48 61
rect 10 8 18 9
rect 34 8 42 9
rect 9 2 19 8
rect 33 2 43 8
rect 10 1 18 2
rect 34 1 42 2
<< labels >>
rlabel metal2 s 12 66 22 74 6 A
port 1 nsew signal input
rlabel metal1 s 12 67 22 73 6 A
port 1 nsew signal input
rlabel metal2 s 38 53 48 61 6 B
port 2 nsew signal input
rlabel metal1 s 38 54 48 60 6 B
port 2 nsew signal input
rlabel metal2 s 10 147 18 155 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 9 148 19 154 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 34 147 42 155 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 33 148 43 154 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 11 106 16 159 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 45 106 50 159 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal1 s 0 147 62 159 6 VDD
port 3 nsew power bidirectional abutment
rlabel metal2 s 10 1 18 9 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 9 2 19 8 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 34 1 42 9 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 33 2 43 8 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 42 -3 47 33 6 VSS
port 4 nsew ground bidirectional
rlabel metal1 s 0 -3 62 9 6 VSS
port 4 nsew ground bidirectional
rlabel metal2 s 26 79 36 87 6 Y
port 5 nsew signal output
rlabel metal1 s 14 16 19 40 6 Y
port 5 nsew signal output
rlabel metal1 s 14 35 33 40 6 Y
port 5 nsew signal output
rlabel metal1 s 28 35 33 140 6 Y
port 5 nsew signal output
rlabel metal1 s 26 80 36 86 6 Y
port 5 nsew signal output
<< properties >>
string FIXED_BBOX 0 -3 62 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
