magic
tech gf180mcuB
timestamp 1667403371
<< metal1 >>
rect 0 111 78 123
rect 28 70 33 111
rect 45 76 50 104
rect 43 70 53 76
rect 62 70 67 111
rect 21 44 31 50
rect 28 12 33 36
rect 45 19 50 70
rect 62 12 67 36
rect 0 0 78 12
<< obsm1 >>
rect 11 65 16 104
rect 11 59 40 65
rect 11 19 16 59
<< metal2 >>
rect 10 118 18 119
rect 34 118 42 119
rect 58 118 66 119
rect 9 112 19 118
rect 33 112 43 118
rect 57 112 67 118
rect 10 111 18 112
rect 34 111 42 112
rect 58 111 66 112
rect 43 69 53 77
rect 22 50 30 51
rect 21 44 31 50
rect 22 43 30 44
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
<< labels >>
rlabel metal2 s 22 43 30 51 6 A
port 1 nsew signal input
rlabel metal2 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal1 s 21 44 31 50 6 A
port 1 nsew signal input
rlabel metal2 s 10 111 18 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 9 112 19 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 34 111 42 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 33 112 43 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 58 111 66 119 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 57 112 67 118 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 28 70 33 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 62 70 67 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal1 s 0 111 78 123 6 VDD
port 2 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 62 0 67 36 6 VSS
port 3 nsew ground bidirectional
rlabel metal1 s 0 0 78 12 6 VSS
port 3 nsew ground bidirectional
rlabel metal2 s 43 69 53 77 6 Y
port 4 nsew signal output
rlabel metal1 s 45 19 50 104 6 Y
port 4 nsew signal output
rlabel metal1 s 43 70 53 76 6 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 78 123
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
