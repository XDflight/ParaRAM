magic
tech gf180mcuB
timestamp 1666464484
<< properties >>
string GDS_END 3127770
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_io/gds/gf180mcu_fd_io.gds
string GDS_START 3124566
<< end >>
