magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -1 7111 1406 7382
rect -1 2294 1525 7111
<< mvnsubdiff >>
rect 751 2649 1023 2668
rect 751 2603 770 2649
rect 1004 2603 1023 2649
rect 751 2584 1023 2603
<< mvnsubdiffcont >>
rect 770 2603 1004 2649
<< polysilicon >>
rect 254 2813 374 2953
rect 254 2767 273 2813
rect 319 2767 374 2813
rect 702 2863 822 3043
rect 926 2863 1046 3028
rect 1150 2863 1270 3046
rect 702 2844 1270 2863
rect 702 2798 1100 2844
rect 1240 2798 1270 2844
rect 702 2779 1270 2798
rect 254 2748 374 2767
rect 702 2333 1270 2352
rect 254 2291 374 2310
rect 254 2245 273 2291
rect 319 2245 374 2291
rect 254 2184 374 2245
rect 702 2287 1100 2333
rect 1240 2287 1270 2333
rect 702 2235 1270 2287
rect 702 2184 822 2235
rect 926 2184 1046 2235
rect 1150 2184 1270 2235
rect 255 2155 373 2184
rect 703 2155 821 2184
rect 927 2155 1045 2184
rect 1151 2155 1269 2184
<< polycontact >>
rect 273 2767 319 2813
rect 1100 2798 1240 2844
rect 273 2245 319 2291
rect 1100 2287 1240 2333
<< metal1 >>
rect 262 2813 330 2824
rect 262 2767 273 2813
rect 319 2767 330 2813
rect 262 2309 330 2767
rect 180 2297 330 2309
rect 180 2245 192 2297
rect 244 2291 330 2297
rect 244 2245 273 2291
rect 319 2245 330 2291
rect 180 2226 330 2245
rect 403 2344 449 3003
rect 851 2660 897 3007
rect 1089 2844 1251 2855
rect 1089 2798 1100 2844
rect 1240 2798 1251 2844
rect 1089 2787 1251 2798
rect 759 2649 1015 2660
rect 759 2603 770 2649
rect 1004 2603 1015 2649
rect 759 2592 1015 2603
rect 1186 2344 1232 2787
rect 403 2333 1251 2344
rect 403 2287 1100 2333
rect 1240 2287 1251 2333
rect 403 2276 1251 2287
rect 403 2062 449 2276
rect 612 2144 688 2156
rect 612 2092 624 2144
rect 676 2092 688 2144
rect 612 2020 688 2092
rect 612 1968 624 2020
rect 676 1968 688 2020
rect 612 1896 688 1968
rect 612 1844 624 1896
rect 676 1844 688 1896
rect 612 1832 688 1844
rect 1060 2144 1136 2156
rect 1060 2092 1072 2144
rect 1124 2092 1136 2144
rect 1060 2020 1136 2092
rect 1060 1968 1072 2020
rect 1124 1968 1136 2020
rect 1060 1896 1136 1968
rect 1060 1844 1072 1896
rect 1124 1844 1136 1896
rect 1060 1832 1136 1844
rect 145 248 260 495
rect 817 248 932 495
rect 1265 248 1380 495
rect 144 -1 260 248
rect 816 -1 932 248
rect 1264 -1 1380 248
<< via1 >>
rect 192 2245 244 2297
rect 624 2092 676 2144
rect 624 1968 676 2020
rect 624 1844 676 1896
rect 1072 2092 1124 2144
rect 1072 1968 1124 2020
rect 1072 1844 1124 1896
<< metal2 >>
rect 180 2297 256 2395
rect 180 2245 192 2297
rect 244 2245 256 2297
rect 180 2233 256 2245
rect 612 2144 688 3302
rect 612 2092 624 2144
rect 676 2092 688 2144
rect 612 2020 688 2092
rect 612 1968 624 2020
rect 676 1968 688 2020
rect 612 1896 688 1968
rect 612 1844 624 1896
rect 676 1844 688 1896
rect 612 1832 688 1844
rect 1060 2144 1136 3313
rect 1060 2092 1072 2144
rect 1124 2092 1136 2144
rect 1060 2020 1136 2092
rect 1060 1968 1072 2020
rect 1124 1968 1136 2020
rect 1060 1896 1136 1968
rect 1060 1844 1072 1896
rect 1124 1844 1136 1896
rect 1060 1832 1136 1844
<< metal3 >>
rect 172 5644 1931 7382
use M1_NWELL4310589983236_64x8m81  M1_NWELL4310589983236_64x8m81_0
timestamp 1666464484
transform 1 0 887 0 1 2626
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_0
timestamp 1666464484
transform 1 0 296 0 1 2790
box 0 0 1 1
use M1_POLY24310589983235_64x8m81  M1_POLY24310589983235_64x8m81_1
timestamp 1666464484
transform 1 0 296 0 1 2268
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_0
timestamp 1666464484
transform 1 0 1170 0 1 2821
box 0 0 1 1
use M1_POLY24310589983237_64x8m81  M1_POLY24310589983237_64x8m81_1
timestamp 1666464484
transform 1 0 1170 0 1 2310
box 0 0 1 1
use M2_M14310589983253_64x8m81  M2_M14310589983253_64x8m81_0
timestamp 1666464484
transform 1 0 874 0 1 6580
box -38 -720 38 720
use M2_M14310589983253_64x8m81  M2_M14310589983253_64x8m81_1
timestamp 1666464484
transform 1 0 1322 0 1 6580
box -38 -720 38 720
use M2_M14310589983253_64x8m81  M2_M14310589983253_64x8m81_2
timestamp 1666464484
transform 1 0 202 0 1 6580
box -38 -720 38 720
use M2_M14310589983255_64x8m81  M2_M14310589983255_64x8m81_0
timestamp 1666464484
transform 1 0 1098 0 1 1994
box 0 0 1 1
use M2_M14310589983255_64x8m81  M2_M14310589983255_64x8m81_1
timestamp 1666464484
transform 1 0 650 0 1 1994
box 0 0 1 1
use M2_M14310589983256_64x8m81  M2_M14310589983256_64x8m81_0
timestamp 1666464484
transform 1 0 218 0 1 2271
box 0 0 1 1
use M2_M14310589983257_64x8m81  M2_M14310589983257_64x8m81_0
timestamp 1666464484
transform 1 0 1098 0 1 4302
box -38 -1092 38 1092
use M2_M14310589983257_64x8m81  M2_M14310589983257_64x8m81_1
timestamp 1666464484
transform 1 0 650 0 1 4302
box -38 -1092 38 1092
use M3_M24310589983254_64x8m81  M3_M24310589983254_64x8m81_0
timestamp 1666464484
transform 1 0 202 0 1 6580
box -38 -720 38 720
use M3_M24310589983254_64x8m81  M3_M24310589983254_64x8m81_1
timestamp 1666464484
transform 1 0 1322 0 1 6580
box -38 -720 38 720
use M3_M24310589983254_64x8m81  M3_M24310589983254_64x8m81_2
timestamp 1666464484
transform 1 0 874 0 1 6580
box -38 -720 38 720
use nmos_5p04310589983258_64x8m81  nmos_5p04310589983258_64x8m81_0
timestamp 1666464484
transform 1 0 926 0 1 340
box -88 -44 208 1860
use nmos_5p04310589983258_64x8m81  nmos_5p04310589983258_64x8m81_1
timestamp 1666464484
transform 1 0 702 0 1 340
box -88 -44 208 1860
use nmos_5p04310589983258_64x8m81  nmos_5p04310589983258_64x8m81_2
timestamp 1666464484
transform 1 0 254 0 1 340
box -88 -44 208 1860
use nmos_5p04310589983258_64x8m81  nmos_5p04310589983258_64x8m81_3
timestamp 1666464484
transform 1 0 1150 0 1 340
box -88 -44 208 1860
use pmos_5p04310589983259_64x8m81  pmos_5p04310589983259_64x8m81_0
timestamp 1666464484
transform 1 0 254 0 1 2971
box -208 -120 328 4120
use pmos_5p04310589983259_64x8m81  pmos_5p04310589983259_64x8m81_1
timestamp 1666464484
transform 1 0 702 0 1 2971
box -208 -120 328 4120
use pmos_5p04310589983259_64x8m81  pmos_5p04310589983259_64x8m81_2
timestamp 1666464484
transform 1 0 926 0 1 2971
box -208 -120 328 4120
use pmos_5p04310589983259_64x8m81  pmos_5p04310589983259_64x8m81_3
timestamp 1666464484
transform 1 0 1150 0 1 2971
box -208 -120 328 4120
<< properties >>
string GDS_END 684794
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 681542
string path 4.370 15.035 4.370 13.055 
<< end >>
