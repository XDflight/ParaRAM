magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 552 312
<< mvpmos >>
rect 0 0 120 192
rect 224 0 344 192
<< mvpdiff >>
rect -88 179 0 192
rect -88 133 -75 179
rect -29 133 0 179
rect -88 59 0 133
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 179 224 192
rect 120 133 149 179
rect 195 133 224 179
rect 120 59 224 133
rect 120 13 149 59
rect 195 13 224 59
rect 120 0 224 13
rect 344 179 432 192
rect 344 133 373 179
rect 419 133 432 179
rect 344 59 432 133
rect 344 13 373 59
rect 419 13 432 59
rect 344 0 432 13
<< mvpdiffc >>
rect -75 133 -29 179
rect -75 13 -29 59
rect 149 133 195 179
rect 149 13 195 59
rect 373 133 419 179
rect 373 13 419 59
<< polysilicon >>
rect 0 192 120 236
rect 224 192 344 236
rect 0 -44 120 0
rect 224 -44 344 0
<< metal1 >>
rect -75 179 -29 192
rect -75 59 -29 133
rect -75 0 -29 13
rect 149 179 195 192
rect 149 59 195 133
rect 149 0 195 13
rect 373 179 419 192
rect 373 59 419 133
rect 373 0 419 13
<< labels >>
flabel metal1 s -52 96 -52 96 0 FreeSans 400 0 0 0 S
flabel metal1 s 396 96 396 96 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 96 172 96 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 164294
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 162568
<< end >>
