magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -208 -120 328 4120
<< mvpmos >>
rect 0 0 120 4000
<< mvpdiff >>
rect -88 3987 0 4000
rect -88 13 -75 3987
rect -29 13 0 3987
rect -88 0 0 13
rect 120 3987 208 4000
rect 120 13 149 3987
rect 195 13 208 3987
rect 120 0 208 13
<< mvpdiffc >>
rect -75 13 -29 3987
rect 149 13 195 3987
<< polysilicon >>
rect 0 4000 120 4044
rect 0 -44 120 0
<< metal1 >>
rect -75 3987 -29 4000
rect -75 0 -29 13
rect 149 3987 195 4000
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 2000 -52 2000 0 FreeSans 400 0 0 0 S
flabel metal1 s 172 2000 172 2000 0 FreeSans 400 0 0 0 D
<< properties >>
string GDS_END 389300
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 383220
<< end >>
