magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -1856 137 1857 175
rect -1856 81 -1820 137
rect -1764 81 -1609 137
rect -1553 81 -1399 137
rect -1343 81 -1188 137
rect -1132 81 -977 137
rect -921 81 -766 137
rect -710 81 -555 137
rect -499 81 -345 137
rect -289 81 -134 137
rect -78 81 78 137
rect 134 81 289 137
rect 345 81 499 137
rect 555 81 710 137
rect 766 81 921 137
rect 977 81 1132 137
rect 1188 81 1343 137
rect 1399 81 1553 137
rect 1609 81 1764 137
rect 1820 81 1857 137
rect -1856 -81 1857 81
rect -1856 -137 -1820 -81
rect -1764 -137 -1609 -81
rect -1553 -137 -1399 -81
rect -1343 -137 -1188 -81
rect -1132 -137 -977 -81
rect -921 -137 -766 -81
rect -710 -137 -555 -81
rect -499 -137 -345 -81
rect -289 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 289 -81
rect 345 -137 499 -81
rect 555 -137 710 -81
rect 766 -137 921 -81
rect 977 -137 1132 -81
rect 1188 -137 1343 -81
rect 1399 -137 1553 -81
rect 1609 -137 1764 -81
rect 1820 -137 1857 -81
rect -1856 -176 1857 -137
<< via2 >>
rect -1820 81 -1764 137
rect -1609 81 -1553 137
rect -1399 81 -1343 137
rect -1188 81 -1132 137
rect -977 81 -921 137
rect -766 81 -710 137
rect -555 81 -499 137
rect -345 81 -289 137
rect -134 81 -78 137
rect 78 81 134 137
rect 289 81 345 137
rect 499 81 555 137
rect 710 81 766 137
rect 921 81 977 137
rect 1132 81 1188 137
rect 1343 81 1399 137
rect 1553 81 1609 137
rect 1764 81 1820 137
rect -1820 -137 -1764 -81
rect -1609 -137 -1553 -81
rect -1399 -137 -1343 -81
rect -1188 -137 -1132 -81
rect -977 -137 -921 -81
rect -766 -137 -710 -81
rect -555 -137 -499 -81
rect -345 -137 -289 -81
rect -134 -137 -78 -81
rect 78 -137 134 -81
rect 289 -137 345 -81
rect 499 -137 555 -81
rect 710 -137 766 -81
rect 921 -137 977 -81
rect 1132 -137 1188 -81
rect 1343 -137 1399 -81
rect 1553 -137 1609 -81
rect 1764 -137 1820 -81
<< metal3 >>
rect -1857 137 1857 176
rect -1857 81 -1820 137
rect -1764 81 -1609 137
rect -1553 81 -1399 137
rect -1343 81 -1188 137
rect -1132 81 -977 137
rect -921 81 -766 137
rect -710 81 -555 137
rect -499 81 -345 137
rect -289 81 -134 137
rect -78 81 78 137
rect 134 81 289 137
rect 345 81 499 137
rect 555 81 710 137
rect 766 81 921 137
rect 977 81 1132 137
rect 1188 81 1343 137
rect 1399 81 1553 137
rect 1609 81 1764 137
rect 1820 81 1857 137
rect -1857 -81 1857 81
rect -1857 -137 -1820 -81
rect -1764 -137 -1609 -81
rect -1553 -137 -1399 -81
rect -1343 -137 -1188 -81
rect -1132 -137 -977 -81
rect -921 -137 -766 -81
rect -710 -137 -555 -81
rect -499 -137 -345 -81
rect -289 -137 -134 -81
rect -78 -137 78 -81
rect 134 -137 289 -81
rect 345 -137 499 -81
rect 555 -137 710 -81
rect 766 -137 921 -81
rect 977 -137 1132 -81
rect 1188 -137 1343 -81
rect 1399 -137 1553 -81
rect 1609 -137 1764 -81
rect 1820 -137 1857 -81
rect -1857 -176 1857 -137
<< properties >>
string GDS_END 951174
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 948738
<< end >>
