magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -1327 -717 1327 717
<< nsubdiff >>
rect -1185 513 1185 570
rect -1185 467 -1130 513
rect -1084 467 -972 513
rect -926 467 -814 513
rect -768 467 -656 513
rect -610 467 -497 513
rect -451 467 -339 513
rect -293 467 -181 513
rect -135 467 -23 513
rect 23 467 135 513
rect 181 467 293 513
rect 339 467 451 513
rect 497 467 610 513
rect 656 467 768 513
rect 814 467 926 513
rect 972 467 1084 513
rect 1130 467 1185 513
rect -1185 350 1185 467
rect -1185 304 -1130 350
rect -1084 304 -972 350
rect -926 304 -814 350
rect -768 304 -656 350
rect -610 304 -497 350
rect -451 304 -339 350
rect -293 304 -181 350
rect -135 304 -23 350
rect 23 304 135 350
rect 181 304 293 350
rect 339 304 451 350
rect 497 304 610 350
rect 656 304 768 350
rect 814 304 926 350
rect 972 304 1084 350
rect 1130 304 1185 350
rect -1185 186 1185 304
rect -1185 140 -1130 186
rect -1084 140 -972 186
rect -926 140 -814 186
rect -768 140 -656 186
rect -610 140 -497 186
rect -451 140 -339 186
rect -293 140 -181 186
rect -135 140 -23 186
rect 23 140 135 186
rect 181 140 293 186
rect 339 140 451 186
rect 497 140 610 186
rect 656 140 768 186
rect 814 140 926 186
rect 972 140 1084 186
rect 1130 140 1185 186
rect -1185 23 1185 140
rect -1185 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1185 23
rect -1185 -140 1185 -23
rect -1185 -186 -1130 -140
rect -1084 -186 -972 -140
rect -926 -186 -814 -140
rect -768 -186 -656 -140
rect -610 -186 -497 -140
rect -451 -186 -339 -140
rect -293 -186 -181 -140
rect -135 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1185 -140
rect -1185 -304 1185 -186
rect -1185 -350 -1130 -304
rect -1084 -350 -972 -304
rect -926 -350 -814 -304
rect -768 -350 -656 -304
rect -610 -350 -497 -304
rect -451 -350 -339 -304
rect -293 -350 -181 -304
rect -135 -350 -23 -304
rect 23 -350 135 -304
rect 181 -350 293 -304
rect 339 -350 451 -304
rect 497 -350 610 -304
rect 656 -350 768 -304
rect 814 -350 926 -304
rect 972 -350 1084 -304
rect 1130 -350 1185 -304
rect -1185 -467 1185 -350
rect -1185 -513 -1130 -467
rect -1084 -513 -972 -467
rect -926 -513 -814 -467
rect -768 -513 -656 -467
rect -610 -513 -497 -467
rect -451 -513 -339 -467
rect -293 -513 -181 -467
rect -135 -513 -23 -467
rect 23 -513 135 -467
rect 181 -513 293 -467
rect 339 -513 451 -467
rect 497 -513 610 -467
rect 656 -513 768 -467
rect 814 -513 926 -467
rect 972 -513 1084 -467
rect 1130 -513 1185 -467
rect -1185 -570 1185 -513
<< nsubdiffcont >>
rect -1130 467 -1084 513
rect -972 467 -926 513
rect -814 467 -768 513
rect -656 467 -610 513
rect -497 467 -451 513
rect -339 467 -293 513
rect -181 467 -135 513
rect -23 467 23 513
rect 135 467 181 513
rect 293 467 339 513
rect 451 467 497 513
rect 610 467 656 513
rect 768 467 814 513
rect 926 467 972 513
rect 1084 467 1130 513
rect -1130 304 -1084 350
rect -972 304 -926 350
rect -814 304 -768 350
rect -656 304 -610 350
rect -497 304 -451 350
rect -339 304 -293 350
rect -181 304 -135 350
rect -23 304 23 350
rect 135 304 181 350
rect 293 304 339 350
rect 451 304 497 350
rect 610 304 656 350
rect 768 304 814 350
rect 926 304 972 350
rect 1084 304 1130 350
rect -1130 140 -1084 186
rect -972 140 -926 186
rect -814 140 -768 186
rect -656 140 -610 186
rect -497 140 -451 186
rect -339 140 -293 186
rect -181 140 -135 186
rect -23 140 23 186
rect 135 140 181 186
rect 293 140 339 186
rect 451 140 497 186
rect 610 140 656 186
rect 768 140 814 186
rect 926 140 972 186
rect 1084 140 1130 186
rect -1130 -23 -1084 23
rect -972 -23 -926 23
rect -814 -23 -768 23
rect -656 -23 -610 23
rect -497 -23 -451 23
rect -339 -23 -293 23
rect -181 -23 -135 23
rect -23 -23 23 23
rect 135 -23 181 23
rect 293 -23 339 23
rect 451 -23 497 23
rect 610 -23 656 23
rect 768 -23 814 23
rect 926 -23 972 23
rect 1084 -23 1130 23
rect -1130 -186 -1084 -140
rect -972 -186 -926 -140
rect -814 -186 -768 -140
rect -656 -186 -610 -140
rect -497 -186 -451 -140
rect -339 -186 -293 -140
rect -181 -186 -135 -140
rect -23 -186 23 -140
rect 135 -186 181 -140
rect 293 -186 339 -140
rect 451 -186 497 -140
rect 610 -186 656 -140
rect 768 -186 814 -140
rect 926 -186 972 -140
rect 1084 -186 1130 -140
rect -1130 -350 -1084 -304
rect -972 -350 -926 -304
rect -814 -350 -768 -304
rect -656 -350 -610 -304
rect -497 -350 -451 -304
rect -339 -350 -293 -304
rect -181 -350 -135 -304
rect -23 -350 23 -304
rect 135 -350 181 -304
rect 293 -350 339 -304
rect 451 -350 497 -304
rect 610 -350 656 -304
rect 768 -350 814 -304
rect 926 -350 972 -304
rect 1084 -350 1130 -304
rect -1130 -513 -1084 -467
rect -972 -513 -926 -467
rect -814 -513 -768 -467
rect -656 -513 -610 -467
rect -497 -513 -451 -467
rect -339 -513 -293 -467
rect -181 -513 -135 -467
rect -23 -513 23 -467
rect 135 -513 181 -467
rect 293 -513 339 -467
rect 451 -513 497 -467
rect 610 -513 656 -467
rect 768 -513 814 -467
rect 926 -513 972 -467
rect 1084 -513 1130 -467
<< metal1 >>
rect -1165 513 1165 550
rect -1165 467 -1130 513
rect -1084 467 -972 513
rect -926 467 -814 513
rect -768 467 -656 513
rect -610 467 -497 513
rect -451 467 -339 513
rect -293 467 -181 513
rect -135 467 -23 513
rect 23 467 135 513
rect 181 467 293 513
rect 339 467 451 513
rect 497 467 610 513
rect 656 467 768 513
rect 814 467 926 513
rect 972 467 1084 513
rect 1130 467 1165 513
rect -1165 350 1165 467
rect -1165 304 -1130 350
rect -1084 304 -972 350
rect -926 304 -814 350
rect -768 304 -656 350
rect -610 304 -497 350
rect -451 304 -339 350
rect -293 304 -181 350
rect -135 304 -23 350
rect 23 304 135 350
rect 181 304 293 350
rect 339 304 451 350
rect 497 304 610 350
rect 656 304 768 350
rect 814 304 926 350
rect 972 304 1084 350
rect 1130 304 1165 350
rect -1165 186 1165 304
rect -1165 140 -1130 186
rect -1084 140 -972 186
rect -926 140 -814 186
rect -768 140 -656 186
rect -610 140 -497 186
rect -451 140 -339 186
rect -293 140 -181 186
rect -135 140 -23 186
rect 23 140 135 186
rect 181 140 293 186
rect 339 140 451 186
rect 497 140 610 186
rect 656 140 768 186
rect 814 140 926 186
rect 972 140 1084 186
rect 1130 140 1165 186
rect -1165 23 1165 140
rect -1165 -23 -1130 23
rect -1084 -23 -972 23
rect -926 -23 -814 23
rect -768 -23 -656 23
rect -610 -23 -497 23
rect -451 -23 -339 23
rect -293 -23 -181 23
rect -135 -23 -23 23
rect 23 -23 135 23
rect 181 -23 293 23
rect 339 -23 451 23
rect 497 -23 610 23
rect 656 -23 768 23
rect 814 -23 926 23
rect 972 -23 1084 23
rect 1130 -23 1165 23
rect -1165 -140 1165 -23
rect -1165 -186 -1130 -140
rect -1084 -186 -972 -140
rect -926 -186 -814 -140
rect -768 -186 -656 -140
rect -610 -186 -497 -140
rect -451 -186 -339 -140
rect -293 -186 -181 -140
rect -135 -186 -23 -140
rect 23 -186 135 -140
rect 181 -186 293 -140
rect 339 -186 451 -140
rect 497 -186 610 -140
rect 656 -186 768 -140
rect 814 -186 926 -140
rect 972 -186 1084 -140
rect 1130 -186 1165 -140
rect -1165 -304 1165 -186
rect -1165 -350 -1130 -304
rect -1084 -350 -972 -304
rect -926 -350 -814 -304
rect -768 -350 -656 -304
rect -610 -350 -497 -304
rect -451 -350 -339 -304
rect -293 -350 -181 -304
rect -135 -350 -23 -304
rect 23 -350 135 -304
rect 181 -350 293 -304
rect 339 -350 451 -304
rect 497 -350 610 -304
rect 656 -350 768 -304
rect 814 -350 926 -304
rect 972 -350 1084 -304
rect 1130 -350 1165 -304
rect -1165 -467 1165 -350
rect -1165 -513 -1130 -467
rect -1084 -513 -972 -467
rect -926 -513 -814 -467
rect -768 -513 -656 -467
rect -610 -513 -497 -467
rect -451 -513 -339 -467
rect -293 -513 -181 -467
rect -135 -513 -23 -467
rect 23 -513 135 -467
rect 181 -513 293 -467
rect 339 -513 451 -467
rect 497 -513 610 -467
rect 656 -513 768 -467
rect 814 -513 926 -467
rect 972 -513 1084 -467
rect 1130 -513 1165 -467
rect -1165 -550 1165 -513
<< properties >>
string GDS_END 661848
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 654868
<< end >>
