magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 1318
<< mvndiff >>
rect -88 1305 0 1318
rect -88 1259 -75 1305
rect -29 1259 0 1305
rect -88 1202 0 1259
rect -88 1156 -75 1202
rect -29 1156 0 1202
rect -88 1099 0 1156
rect -88 1053 -75 1099
rect -29 1053 0 1099
rect -88 995 0 1053
rect -88 949 -75 995
rect -29 949 0 995
rect -88 891 0 949
rect -88 845 -75 891
rect -29 845 0 891
rect -88 787 0 845
rect -88 741 -75 787
rect -29 741 0 787
rect -88 683 0 741
rect -88 637 -75 683
rect -29 637 0 683
rect -88 579 0 637
rect -88 533 -75 579
rect -29 533 0 579
rect -88 475 0 533
rect -88 429 -75 475
rect -29 429 0 475
rect -88 371 0 429
rect -88 325 -75 371
rect -29 325 0 371
rect -88 267 0 325
rect -88 221 -75 267
rect -29 221 0 267
rect -88 163 0 221
rect -88 117 -75 163
rect -29 117 0 163
rect -88 59 0 117
rect -88 13 -75 59
rect -29 13 0 59
rect -88 0 0 13
rect 120 1305 208 1318
rect 120 1259 149 1305
rect 195 1259 208 1305
rect 120 1202 208 1259
rect 120 1156 149 1202
rect 195 1156 208 1202
rect 120 1099 208 1156
rect 120 1053 149 1099
rect 195 1053 208 1099
rect 120 995 208 1053
rect 120 949 149 995
rect 195 949 208 995
rect 120 891 208 949
rect 120 845 149 891
rect 195 845 208 891
rect 120 787 208 845
rect 120 741 149 787
rect 195 741 208 787
rect 120 683 208 741
rect 120 637 149 683
rect 195 637 208 683
rect 120 579 208 637
rect 120 533 149 579
rect 195 533 208 579
rect 120 475 208 533
rect 120 429 149 475
rect 195 429 208 475
rect 120 371 208 429
rect 120 325 149 371
rect 195 325 208 371
rect 120 267 208 325
rect 120 221 149 267
rect 195 221 208 267
rect 120 163 208 221
rect 120 117 149 163
rect 195 117 208 163
rect 120 59 208 117
rect 120 13 149 59
rect 195 13 208 59
rect 120 0 208 13
<< mvndiffc >>
rect -75 1259 -29 1305
rect -75 1156 -29 1202
rect -75 1053 -29 1099
rect -75 949 -29 995
rect -75 845 -29 891
rect -75 741 -29 787
rect -75 637 -29 683
rect -75 533 -29 579
rect -75 429 -29 475
rect -75 325 -29 371
rect -75 221 -29 267
rect -75 117 -29 163
rect -75 13 -29 59
rect 149 1259 195 1305
rect 149 1156 195 1202
rect 149 1053 195 1099
rect 149 949 195 995
rect 149 845 195 891
rect 149 741 195 787
rect 149 637 195 683
rect 149 533 195 579
rect 149 429 195 475
rect 149 325 195 371
rect 149 221 195 267
rect 149 117 195 163
rect 149 13 195 59
<< polysilicon >>
rect 0 1318 120 1362
rect 0 -44 120 0
<< metal1 >>
rect -75 1305 -29 1318
rect -75 1202 -29 1259
rect -75 1099 -29 1156
rect -75 995 -29 1053
rect -75 891 -29 949
rect -75 787 -29 845
rect -75 683 -29 741
rect -75 579 -29 637
rect -75 475 -29 533
rect -75 371 -29 429
rect -75 267 -29 325
rect -75 163 -29 221
rect -75 59 -29 117
rect -75 0 -29 13
rect 149 1305 195 1318
rect 149 1202 195 1259
rect 149 1099 195 1156
rect 149 995 195 1053
rect 149 891 195 949
rect 149 787 195 845
rect 149 683 195 741
rect 149 579 195 637
rect 149 475 195 533
rect 149 371 195 429
rect 149 267 195 325
rect 149 163 195 221
rect 149 59 195 117
rect 149 0 195 13
<< labels >>
flabel metal1 s -52 659 -52 659 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 659 172 659 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 645520
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 642960
<< end >>
