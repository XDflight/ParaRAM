magic
tech gf180mcuA
timestamp 1667403424
<< metal1 >>
rect 0 150 280 162
rect 28 109 33 150
rect 30 83 40 89
rect 12 70 22 76
rect 96 109 101 150
rect 130 109 135 150
rect 72 83 125 89
rect 92 70 102 76
rect 215 109 220 150
rect 232 89 237 143
rect 247 109 252 150
rect 191 83 201 89
rect 232 83 240 89
rect 174 70 184 76
rect 47 57 57 63
rect 28 12 33 36
rect 133 44 143 50
rect 96 12 101 36
rect 130 12 135 29
rect 201 44 211 50
rect 215 12 220 36
rect 232 19 237 83
rect 264 64 269 143
rect 264 63 272 64
rect 264 57 275 63
rect 264 56 272 57
rect 247 12 252 36
rect 264 19 269 56
rect 0 0 280 12
<< obsm1 >>
rect 11 104 16 143
rect 45 104 50 143
rect 11 99 50 104
rect 62 63 67 143
rect 113 104 118 143
rect 147 104 152 143
rect 113 99 152 104
rect 164 63 169 143
rect 62 57 159 63
rect 164 57 227 63
rect 11 41 50 46
rect 11 19 16 41
rect 45 19 50 41
rect 62 19 67 57
rect 113 34 152 39
rect 113 19 118 34
rect 147 19 152 34
rect 164 19 169 57
rect 249 57 259 63
<< metal2 >>
rect 10 157 18 158
rect 34 157 42 158
rect 58 157 66 158
rect 82 157 90 158
rect 106 157 114 158
rect 130 157 138 158
rect 154 157 162 158
rect 178 157 186 158
rect 202 157 210 158
rect 226 157 234 158
rect 250 157 258 158
rect 9 151 19 157
rect 33 151 43 157
rect 57 151 67 157
rect 81 151 91 157
rect 105 151 115 157
rect 129 151 139 157
rect 153 151 163 157
rect 177 151 187 157
rect 201 151 211 157
rect 225 151 235 157
rect 249 151 259 157
rect 10 150 18 151
rect 34 150 42 151
rect 58 150 66 151
rect 82 150 90 151
rect 106 150 114 151
rect 130 150 138 151
rect 154 150 162 151
rect 178 150 186 151
rect 202 150 210 151
rect 226 150 234 151
rect 250 150 258 151
rect 31 89 39 90
rect 73 89 81 90
rect 116 89 124 90
rect 192 89 200 90
rect 231 89 239 90
rect 30 83 82 89
rect 115 83 201 89
rect 230 83 240 89
rect 31 82 39 83
rect 73 82 81 83
rect 116 82 124 83
rect 192 82 200 83
rect 231 82 239 83
rect 13 76 21 77
rect 93 76 101 77
rect 175 76 183 77
rect 12 70 184 76
rect 13 69 21 70
rect 93 69 101 70
rect 175 69 183 70
rect 48 63 56 64
rect 266 63 274 64
rect 47 57 57 63
rect 265 57 275 63
rect 48 56 56 57
rect 266 56 274 57
rect 49 50 55 56
rect 134 50 142 51
rect 202 50 210 51
rect 49 44 211 50
rect 134 43 142 44
rect 202 43 210 44
rect 135 42 141 43
rect 203 42 209 43
rect 10 11 18 12
rect 34 11 42 12
rect 58 11 66 12
rect 82 11 90 12
rect 106 11 114 12
rect 130 11 138 12
rect 154 11 162 12
rect 178 11 186 12
rect 202 11 210 12
rect 226 11 234 12
rect 250 11 258 12
rect 9 5 19 11
rect 33 5 43 11
rect 57 5 67 11
rect 81 5 91 11
rect 105 5 115 11
rect 129 5 139 11
rect 153 5 163 11
rect 177 5 187 11
rect 201 5 211 11
rect 225 5 235 11
rect 249 5 259 11
rect 10 4 18 5
rect 34 4 42 5
rect 58 4 66 5
rect 82 4 90 5
rect 106 4 114 5
rect 130 4 138 5
rect 154 4 162 5
rect 178 4 186 5
rect 202 4 210 5
rect 226 4 234 5
rect 250 4 258 5
<< obsm2 >>
rect 150 63 158 64
rect 250 63 258 64
rect 149 57 259 63
rect 150 56 158 57
rect 250 56 258 57
rect 251 55 257 56
<< labels >>
rlabel metal2 s 13 69 21 77 6 A
port 1 nsew signal input
rlabel metal2 s 93 69 101 77 6 A
port 1 nsew signal input
rlabel metal2 s 175 69 183 77 6 A
port 1 nsew signal input
rlabel metal2 s 12 70 184 76 6 A
port 1 nsew signal input
rlabel metal1 s 12 70 22 76 6 A
port 1 nsew signal input
rlabel metal1 s 92 70 102 76 6 A
port 1 nsew signal input
rlabel metal1 s 174 70 184 76 6 A
port 1 nsew signal input
rlabel metal2 s 31 82 39 90 6 B
port 2 nsew signal input
rlabel metal2 s 73 82 81 90 6 B
port 2 nsew signal input
rlabel metal2 s 30 83 82 89 6 B
port 2 nsew signal input
rlabel metal2 s 116 82 124 90 6 B
port 2 nsew signal input
rlabel metal2 s 192 82 200 90 6 B
port 2 nsew signal input
rlabel metal2 s 115 83 201 89 6 B
port 2 nsew signal input
rlabel metal1 s 30 83 40 89 6 B
port 2 nsew signal input
rlabel metal1 s 72 83 125 89 6 B
port 2 nsew signal input
rlabel metal1 s 191 83 201 89 6 B
port 2 nsew signal input
rlabel metal2 s 49 44 55 64 6 CI
port 3 nsew signal input
rlabel metal2 s 48 56 56 64 6 CI
port 3 nsew signal input
rlabel metal2 s 47 57 57 63 6 CI
port 3 nsew signal input
rlabel metal2 s 135 42 141 51 6 CI
port 3 nsew signal input
rlabel metal2 s 134 43 142 51 6 CI
port 3 nsew signal input
rlabel metal2 s 203 42 209 51 6 CI
port 3 nsew signal input
rlabel metal2 s 202 43 210 51 6 CI
port 3 nsew signal input
rlabel metal2 s 49 44 211 50 6 CI
port 3 nsew signal input
rlabel metal1 s 47 57 57 63 6 CI
port 3 nsew signal input
rlabel metal1 s 133 44 143 50 6 CI
port 3 nsew signal input
rlabel metal1 s 201 44 211 50 6 CI
port 3 nsew signal input
rlabel metal2 s 266 56 274 64 6 CO
port 4 nsew signal output
rlabel metal2 s 265 57 275 63 6 CO
port 4 nsew signal output
rlabel metal1 s 264 19 269 143 6 CO
port 4 nsew signal output
rlabel metal1 s 264 56 272 64 6 CO
port 4 nsew signal output
rlabel metal1 s 264 57 275 63 6 CO
port 4 nsew signal output
rlabel metal2 s 231 82 239 90 6 S
port 5 nsew signal output
rlabel metal2 s 230 83 240 89 6 S
port 5 nsew signal output
rlabel metal1 s 232 19 237 143 6 S
port 5 nsew signal output
rlabel metal1 s 232 83 240 89 6 S
port 5 nsew signal output
rlabel metal2 s 10 150 18 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 9 151 19 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 34 150 42 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 33 151 43 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 58 150 66 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 57 151 67 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 82 150 90 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 81 151 91 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 106 150 114 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 105 151 115 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 130 150 138 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 129 151 139 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 154 150 162 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 153 151 163 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 178 150 186 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 177 151 187 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 202 150 210 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 201 151 211 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 226 150 234 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 225 151 235 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 250 150 258 158 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 249 151 259 157 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 28 109 33 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 96 109 101 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 130 109 135 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 215 109 220 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 247 109 252 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal1 s 0 150 280 162 6 VDD
port 6 nsew power bidirectional abutment
rlabel metal2 s 10 4 18 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 9 5 19 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 34 4 42 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 33 5 43 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 58 4 66 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 57 5 67 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 82 4 90 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 81 5 91 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 106 4 114 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 105 5 115 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 130 4 138 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 129 5 139 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 154 4 162 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 153 5 163 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 178 4 186 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 177 5 187 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 202 4 210 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 201 5 211 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 226 4 234 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 225 5 235 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 250 4 258 12 6 VSS
port 7 nsew ground bidirectional
rlabel metal2 s 249 5 259 11 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 28 0 33 36 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 96 0 101 36 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 130 0 135 29 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 215 0 220 36 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 247 0 252 36 6 VSS
port 7 nsew ground bidirectional
rlabel metal1 s 0 0 280 12 6 VSS
port 7 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 280 162
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
