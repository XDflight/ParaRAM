magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 2016 844
rect 69 506 115 724
rect 174 472 855 536
rect 174 353 242 472
rect 319 360 700 424
rect 786 365 855 472
rect 993 506 1039 724
rect 1217 536 1263 678
rect 1421 587 1467 724
rect 1635 536 1681 678
rect 1849 588 1895 724
rect 1217 472 1892 536
rect 1841 308 1892 472
rect 49 60 95 214
rect 497 60 543 214
rect 1197 253 1892 308
rect 1197 252 1691 253
rect 945 60 991 214
rect 1197 106 1243 252
rect 1421 60 1467 197
rect 1645 106 1691 252
rect 1869 60 1915 196
rect 0 -60 2016 60
<< obsm1 >>
rect 470 589 947 643
rect 901 419 947 589
rect 901 365 1792 419
rect 901 314 947 365
rect 273 265 947 314
rect 273 106 319 265
rect 721 106 767 265
<< labels >>
rlabel metal1 s 319 360 700 424 6 A1
port 1 nsew default input
rlabel metal1 s 174 472 855 536 6 A2
port 2 nsew default input
rlabel metal1 s 786 365 855 472 6 A2
port 2 nsew default input
rlabel metal1 s 174 365 242 472 6 A2
port 2 nsew default input
rlabel metal1 s 174 353 242 365 6 A2
port 2 nsew default input
rlabel metal1 s 1635 536 1681 678 6 Z
port 3 nsew default output
rlabel metal1 s 1217 536 1263 678 6 Z
port 3 nsew default output
rlabel metal1 s 1217 472 1892 536 6 Z
port 3 nsew default output
rlabel metal1 s 1841 308 1892 472 6 Z
port 3 nsew default output
rlabel metal1 s 1197 253 1892 308 6 Z
port 3 nsew default output
rlabel metal1 s 1197 252 1691 253 6 Z
port 3 nsew default output
rlabel metal1 s 1645 106 1691 252 6 Z
port 3 nsew default output
rlabel metal1 s 1197 106 1243 252 6 Z
port 3 nsew default output
rlabel metal1 s 0 724 2016 844 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1849 588 1895 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1421 588 1467 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 993 588 1039 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 69 588 115 724 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 1421 587 1467 588 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 993 587 1039 588 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 69 587 115 588 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 993 506 1039 587 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 69 506 115 587 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 945 197 991 214 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 497 197 543 214 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 49 197 95 214 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1421 196 1467 197 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 945 196 991 197 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 497 196 543 197 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 49 196 95 197 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1869 60 1915 196 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 1421 60 1467 196 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 196 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 196 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 196 6 VSS
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 2016 60 8 VSS
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2016 784
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 151300
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 146738
<< end >>
