magic
tech gf180mcuC
magscale 1 5
timestamp 1667403444
<< checkpaint >>
rect 14000 14000 36500 36500
<< metal3 >>
rect 15000 26374 16500 35500
tri 16500 26374 17122 26996 sw
tri 15000 25610 15764 26374 ne
rect 15764 25610 17122 26374
tri 17122 25610 17886 26374 sw
tri 15764 23488 17886 25610 ne
tri 17886 23488 20008 25610 sw
tri 17886 21366 20008 23488 ne
tri 20008 21366 22130 23488 sw
tri 20008 19244 22130 21366 ne
tri 22130 19244 24252 21366 sw
tri 22130 17122 24252 19244 ne
tri 24252 17122 26374 19244 sw
tri 24252 15000 26374 17122 ne
tri 26374 16500 26996 17122 sw
rect 26374 15000 35500 16500
<< end >>
