magic
tech gf180mcuB
magscale 1 10
timestamp 1667403392
<< checkpaint >>
rect 40800 40800 73000 73000
<< metal4 >>
rect 42800 58097 45800 71000
tri 45800 58097 47053 59350 sw
tri 42800 55559 45338 58097 ne
rect 45338 55559 47053 58097
tri 47053 55559 49591 58097 sw
tri 45338 51306 49591 55559 ne
tri 49591 51306 53844 55559 sw
tri 49591 47053 53844 51306 ne
tri 53844 47053 58097 51306 sw
tri 53844 42800 58097 47053 ne
tri 58097 45799 59351 47053 sw
rect 58097 42800 71000 45799
<< end >>
