magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -653 23 653 42
rect -653 -23 -634 23
rect 634 -23 653 23
rect -653 -42 653 -23
<< psubdiffcont >>
rect -634 -23 634 23
<< metal1 >>
rect -645 23 645 34
rect -645 -23 -634 23
rect 634 -23 645 23
rect -645 -34 645 -23
<< properties >>
string GDS_END 2028686
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 2027594
<< end >>
