magic
tech gf180mcuC
timestamp 1666464484
<< metal1 >>
rect -2 147 94 159
rect 9 106 14 147
rect 9 54 19 60
rect 43 74 48 140
rect 60 100 65 140
rect 58 92 68 100
rect 43 66 55 74
rect 9 9 14 33
rect 43 16 48 66
rect 60 16 65 92
rect 77 87 82 140
rect 73 79 83 87
rect 77 16 82 79
rect -2 -3 94 9
<< obsm1 >>
rect 26 86 31 140
rect 26 80 38 86
rect 26 47 31 80
rect 26 41 38 47
rect 26 16 31 41
<< metal2 >>
rect 8 154 16 155
rect 32 154 40 155
rect 56 154 64 155
rect 7 148 17 154
rect 31 148 41 154
rect 55 148 65 154
rect 8 147 16 148
rect 32 147 40 148
rect 56 147 64 148
rect 58 92 68 100
rect 73 79 83 87
rect 45 66 55 74
rect 9 53 19 61
rect 8 8 16 9
rect 32 8 40 9
rect 56 8 64 9
rect 7 2 17 8
rect 31 2 41 8
rect 55 2 65 8
rect 8 1 16 2
rect 32 1 40 2
rect 56 1 64 2
<< labels >>
rlabel metal2 s 45 66 55 74 6 A
port 1 nsew signal input
rlabel metal1 s 43 16 48 140 6 A
port 1 nsew signal input
rlabel metal1 s 43 66 55 74 6 A
port 1 nsew signal input
rlabel metal2 s 73 79 83 87 6 B
port 2 nsew signal input
rlabel metal1 s 77 16 82 140 6 B
port 2 nsew signal input
rlabel metal1 s 73 79 83 87 6 B
port 2 nsew signal input
rlabel metal2 s 9 53 19 61 6 Sel
port 3 nsew signal output
rlabel metal1 s 9 54 19 60 6 Sel
port 3 nsew signal output
rlabel metal2 s 8 147 16 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 7 148 17 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 32 147 40 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 31 148 41 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 56 147 64 155 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 55 148 65 154 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s 9 106 14 159 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal1 s -2 147 94 159 6 VDD
port 4 nsew power bidirectional abutment
rlabel metal2 s 8 1 16 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 7 2 17 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 32 1 40 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 31 2 41 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 56 1 64 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 55 2 65 8 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s 9 -3 14 33 6 VSS
port 5 nsew ground bidirectional
rlabel metal1 s -2 -3 94 9 6 VSS
port 5 nsew ground bidirectional
rlabel metal2 s 58 92 68 100 6 Y
port 6 nsew signal output
rlabel metal1 s 60 16 65 140 6 Y
port 6 nsew signal output
rlabel metal1 s 58 92 68 100 6 Y
port 6 nsew signal output
<< properties >>
string FIXED_BBOX -2 -3 94 159
string LEFclass CORE
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
<< end >>
