magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 1044 88 1116
rect -31 -74 88 -1
use nmos_5p04310589983269_64x8m81  nmos_5p04310589983269_64x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 208 1088
<< properties >>
string GDS_END 78474
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 78224
<< end >>
