magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -60 -407 2159 1742
<< pmos >>
rect 206 507 994 1606
rect 1106 507 1894 1606
<< pdiff >>
rect 81 1563 206 1606
rect 81 1517 127 1563
rect 173 1517 206 1563
rect 81 1402 206 1517
rect 81 1356 127 1402
rect 173 1356 206 1402
rect 81 1242 206 1356
rect 81 1196 127 1242
rect 173 1196 206 1242
rect 81 1082 206 1196
rect 81 1036 127 1082
rect 173 1036 206 1082
rect 81 921 206 1036
rect 81 875 127 921
rect 173 875 206 921
rect 81 759 206 875
rect 81 713 127 759
rect 173 713 206 759
rect 81 596 206 713
rect 81 550 127 596
rect 173 550 206 596
rect 81 507 206 550
rect 994 1563 1106 1606
rect 994 1517 1027 1563
rect 1073 1517 1106 1563
rect 994 1402 1106 1517
rect 994 1356 1027 1402
rect 1073 1356 1106 1402
rect 994 1242 1106 1356
rect 994 1196 1027 1242
rect 1073 1196 1106 1242
rect 994 1082 1106 1196
rect 994 1036 1027 1082
rect 1073 1036 1106 1082
rect 994 921 1106 1036
rect 994 875 1027 921
rect 1073 875 1106 921
rect 994 759 1106 875
rect 994 713 1027 759
rect 1073 713 1106 759
rect 994 596 1106 713
rect 994 550 1027 596
rect 1073 550 1106 596
rect 994 507 1106 550
rect 1894 1563 2019 1606
rect 1894 1517 1927 1563
rect 1973 1517 2019 1563
rect 1894 1402 2019 1517
rect 1894 1356 1927 1402
rect 1973 1356 2019 1402
rect 1894 1242 2019 1356
rect 1894 1196 1927 1242
rect 1973 1196 2019 1242
rect 1894 1082 2019 1196
rect 1894 1036 1927 1082
rect 1973 1036 2019 1082
rect 1894 921 2019 1036
rect 1894 875 1927 921
rect 1973 875 2019 921
rect 1894 759 2019 875
rect 1894 713 1927 759
rect 1973 713 2019 759
rect 1894 596 2019 713
rect 1894 550 1927 596
rect 1973 550 2019 596
rect 1894 507 2019 550
<< pdiffc >>
rect 127 1517 173 1563
rect 127 1356 173 1402
rect 127 1196 173 1242
rect 127 1036 173 1082
rect 127 875 173 921
rect 127 713 173 759
rect 127 550 173 596
rect 1027 1517 1073 1563
rect 1027 1356 1073 1402
rect 1027 1196 1073 1242
rect 1027 1036 1073 1082
rect 1027 875 1073 921
rect 1027 713 1073 759
rect 1027 550 1073 596
rect 1927 1517 1973 1563
rect 1927 1356 1973 1402
rect 1927 1196 1973 1242
rect 1927 1036 1973 1082
rect 1927 875 1973 921
rect 1927 713 1973 759
rect 1927 550 1973 596
<< psubdiff >>
rect 49 2070 2050 2124
rect 49 2024 211 2070
rect 257 2024 374 2070
rect 420 2024 537 2070
rect 583 2024 700 2070
rect 746 2024 864 2070
rect 910 2024 1027 2070
rect 1073 2024 1190 2070
rect 1236 2024 1354 2070
rect 1400 2024 1517 2070
rect 1563 2024 1680 2070
rect 1726 2024 1843 2070
rect 1889 2024 2050 2070
rect 49 1969 2050 2024
<< nsubdiff >>
rect 83 243 2016 297
rect 83 197 211 243
rect 257 197 374 243
rect 420 197 537 243
rect 583 197 700 243
rect 746 197 864 243
rect 910 197 1027 243
rect 1073 197 1190 243
rect 1236 197 1354 243
rect 1400 197 1517 243
rect 1563 197 1680 243
rect 1726 197 1843 243
rect 1889 197 2016 243
rect 83 78 2016 197
<< psubdiffcont >>
rect 211 2024 257 2070
rect 374 2024 420 2070
rect 537 2024 583 2070
rect 700 2024 746 2070
rect 864 2024 910 2070
rect 1027 2024 1073 2070
rect 1190 2024 1236 2070
rect 1354 2024 1400 2070
rect 1517 2024 1563 2070
rect 1680 2024 1726 2070
rect 1843 2024 1889 2070
<< nsubdiffcont >>
rect 211 197 257 243
rect 374 197 420 243
rect 537 197 583 243
rect 700 197 746 243
rect 864 197 910 243
rect 1027 197 1073 243
rect 1190 197 1236 243
rect 1354 197 1400 243
rect 1517 197 1563 243
rect 1680 197 1726 243
rect 1843 197 1889 243
<< polysilicon >>
rect 206 1764 994 1808
rect 206 1718 333 1764
rect 379 1718 496 1764
rect 542 1718 660 1764
rect 706 1718 823 1764
rect 869 1718 994 1764
rect 206 1606 994 1718
rect 1106 1764 1894 1808
rect 1106 1718 1233 1764
rect 1279 1718 1396 1764
rect 1442 1718 1560 1764
rect 1606 1718 1723 1764
rect 1769 1718 1894 1764
rect 1106 1606 1894 1718
rect 206 436 994 507
rect 1106 436 1894 507
<< polycontact >>
rect 333 1718 379 1764
rect 496 1718 542 1764
rect 660 1718 706 1764
rect 823 1718 869 1764
rect 1233 1718 1279 1764
rect 1396 1718 1442 1764
rect 1560 1718 1606 1764
rect 1723 1718 1769 1764
<< metal1 >>
rect 49 2070 2050 2124
rect 49 2024 211 2070
rect 257 2024 374 2070
rect 420 2024 537 2070
rect 583 2024 700 2070
rect 746 2024 864 2070
rect 910 2035 1027 2070
rect 1073 2035 1190 2070
rect 910 2024 1024 2035
rect 1076 2024 1190 2035
rect 1236 2024 1354 2070
rect 1400 2024 1517 2070
rect 1563 2024 1680 2070
rect 1726 2024 1843 2070
rect 1889 2024 2050 2070
rect 49 1983 1024 2024
rect 1076 1983 2050 2024
rect 49 1824 2050 1983
rect 49 1772 1024 1824
rect 1076 1772 2050 1824
rect 49 1764 2050 1772
rect 49 1718 333 1764
rect 379 1718 496 1764
rect 542 1718 660 1764
rect 706 1718 823 1764
rect 869 1718 1233 1764
rect 1279 1718 1396 1764
rect 1442 1718 1560 1764
rect 1606 1718 1723 1764
rect 1769 1718 2050 1764
rect 49 1684 2050 1718
rect 83 1563 216 1597
rect 83 1517 127 1563
rect 173 1517 216 1563
rect 83 1402 216 1517
rect 83 1356 127 1402
rect 173 1356 216 1402
rect 83 1336 216 1356
rect 983 1563 1116 1597
rect 983 1517 1027 1563
rect 1073 1517 1116 1563
rect 983 1402 1116 1517
rect 983 1356 1027 1402
rect 1073 1356 1116 1402
rect 983 1336 1116 1356
rect 1883 1563 2016 1597
rect 1883 1517 1927 1563
rect 1973 1517 2016 1563
rect 1883 1402 2016 1517
rect 1883 1356 1927 1402
rect 1973 1356 2016 1402
rect 1883 1336 2016 1356
rect 83 1298 217 1336
rect 83 1246 124 1298
rect 176 1246 217 1298
rect 83 1242 217 1246
rect 83 1196 127 1242
rect 173 1196 217 1242
rect 83 1087 217 1196
rect 83 1035 124 1087
rect 176 1035 217 1087
rect 83 921 217 1035
rect 83 875 127 921
rect 173 875 217 921
rect 83 823 124 875
rect 176 823 217 875
rect 83 759 217 823
rect 83 713 127 759
rect 173 713 217 759
rect 83 664 217 713
rect 83 612 124 664
rect 176 612 217 664
rect 83 596 217 612
rect 83 550 127 596
rect 173 574 217 596
rect 983 1298 1117 1336
rect 983 1246 1024 1298
rect 1076 1246 1117 1298
rect 983 1242 1117 1246
rect 983 1196 1027 1242
rect 1073 1196 1117 1242
rect 983 1087 1117 1196
rect 983 1035 1024 1087
rect 1076 1035 1117 1087
rect 983 921 1117 1035
rect 983 875 1027 921
rect 1073 875 1117 921
rect 983 823 1024 875
rect 1076 823 1117 875
rect 983 759 1117 823
rect 983 713 1027 759
rect 1073 713 1117 759
rect 983 664 1117 713
rect 983 612 1024 664
rect 1076 612 1117 664
rect 983 596 1117 612
rect 173 550 216 574
rect 83 515 216 550
rect 983 550 1027 596
rect 1073 574 1117 596
rect 1883 1298 2017 1336
rect 1883 1246 1924 1298
rect 1976 1246 2017 1298
rect 1883 1242 2017 1246
rect 1883 1196 1927 1242
rect 1973 1196 2017 1242
rect 1883 1087 2017 1196
rect 1883 1035 1924 1087
rect 1976 1035 2017 1087
rect 1883 921 2017 1035
rect 1883 875 1927 921
rect 1973 875 2017 921
rect 1883 823 1924 875
rect 1976 823 2017 875
rect 1883 759 2017 823
rect 1883 713 1927 759
rect 1973 713 2017 759
rect 1883 664 2017 713
rect 1883 612 1924 664
rect 1976 612 2017 664
rect 1883 596 2017 612
rect 1073 550 1116 574
rect 983 515 1116 550
rect 1883 550 1927 596
rect 1973 574 2017 596
rect 1973 550 2016 574
rect 1883 515 2016 550
rect 83 243 2016 297
rect 83 197 211 243
rect 257 197 374 243
rect 420 197 537 243
rect 583 197 700 243
rect 746 197 864 243
rect 910 197 1027 243
rect 1073 197 1190 243
rect 1236 197 1354 243
rect 1400 197 1517 243
rect 1563 197 1680 243
rect 1726 197 1843 243
rect 1889 197 2016 243
rect 83 78 2016 197
<< via1 >>
rect 1024 2024 1027 2035
rect 1027 2024 1073 2035
rect 1073 2024 1076 2035
rect 1024 1983 1076 2024
rect 1024 1772 1076 1824
rect 124 1246 176 1298
rect 124 1082 176 1087
rect 124 1036 127 1082
rect 127 1036 173 1082
rect 173 1036 176 1082
rect 124 1035 176 1036
rect 124 823 176 875
rect 124 612 176 664
rect 1024 1246 1076 1298
rect 1024 1082 1076 1087
rect 1024 1036 1027 1082
rect 1027 1036 1073 1082
rect 1073 1036 1076 1082
rect 1024 1035 1076 1036
rect 1024 823 1076 875
rect 1024 612 1076 664
rect 1924 1246 1976 1298
rect 1924 1082 1976 1087
rect 1924 1036 1927 1082
rect 1927 1036 1973 1082
rect 1973 1036 1976 1082
rect 1924 1035 1976 1036
rect 1924 823 1976 875
rect 1924 612 1976 664
<< metal2 >>
rect 983 2035 1117 2074
rect 983 1983 1024 2035
rect 1076 1983 1117 2035
rect 983 1826 1117 1983
rect 983 1770 1022 1826
rect 1078 1770 1117 1826
rect 983 1734 1117 1770
rect 49 1300 2050 1395
rect 49 1244 122 1300
rect 178 1298 1922 1300
rect 178 1246 1024 1298
rect 1076 1246 1922 1298
rect 178 1244 1922 1246
rect 1978 1244 2050 1300
rect 49 1089 2050 1244
rect 49 1033 122 1089
rect 178 1087 1922 1089
rect 178 1035 1024 1087
rect 1076 1035 1922 1087
rect 178 1033 1922 1035
rect 1978 1033 2050 1089
rect 49 877 2050 1033
rect 49 821 122 877
rect 178 875 1922 877
rect 178 823 1024 875
rect 1076 823 1922 875
rect 178 821 1922 823
rect 1978 821 2050 877
rect 49 666 2050 821
rect 49 610 122 666
rect 178 664 1922 666
rect 178 612 1024 664
rect 1076 612 1922 664
rect 178 610 1922 612
rect 1978 610 2050 666
rect 49 515 2050 610
<< via2 >>
rect 1022 1824 1078 1826
rect 1022 1772 1024 1824
rect 1024 1772 1076 1824
rect 1076 1772 1078 1824
rect 1022 1770 1078 1772
rect 122 1298 178 1300
rect 1922 1298 1978 1300
rect 122 1246 124 1298
rect 124 1246 176 1298
rect 176 1246 178 1298
rect 1922 1246 1924 1298
rect 1924 1246 1976 1298
rect 1976 1246 1978 1298
rect 122 1244 178 1246
rect 1922 1244 1978 1246
rect 122 1087 178 1089
rect 1922 1087 1978 1089
rect 122 1035 124 1087
rect 124 1035 176 1087
rect 176 1035 178 1087
rect 1922 1035 1924 1087
rect 1924 1035 1976 1087
rect 1976 1035 1978 1087
rect 122 1033 178 1035
rect 1922 1033 1978 1035
rect 122 875 178 877
rect 1922 875 1978 877
rect 122 823 124 875
rect 124 823 176 875
rect 176 823 178 875
rect 1922 823 1924 875
rect 1924 823 1976 875
rect 1976 823 1978 875
rect 122 821 178 823
rect 1922 821 1978 823
rect 122 664 178 666
rect 1922 664 1978 666
rect 122 612 124 664
rect 124 612 176 664
rect 176 612 178 664
rect 1922 612 1924 664
rect 1924 612 1976 664
rect 1976 612 1978 664
rect 122 610 178 612
rect 1922 610 1978 612
<< metal3 >>
rect 49 1300 250 5567
rect 49 1244 122 1300
rect 178 1244 250 1300
rect 49 1089 250 1244
rect 49 1033 122 1089
rect 178 1033 250 1089
rect 49 877 250 1033
rect 49 821 122 877
rect 178 821 250 877
rect 49 666 250 821
rect 49 610 122 666
rect 178 610 250 666
rect 49 -1 250 610
rect 489 -1 690 5567
rect 949 1826 1150 5567
rect 949 1770 1022 1826
rect 1078 1770 1150 1826
rect 949 -1 1150 1770
rect 1409 -1 1611 5567
rect 1849 1300 2050 5567
rect 1849 1244 1922 1300
rect 1978 1244 2050 1300
rect 1849 1089 2050 1244
rect 1849 1033 1922 1089
rect 1978 1033 2050 1089
rect 1849 877 2050 1033
rect 1849 821 1922 877
rect 1978 821 2050 877
rect 1849 666 2050 821
rect 1849 610 1922 666
rect 1978 610 2050 666
rect 1849 -1 2050 610
<< properties >>
string GDS_END 1328804
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 1321248
<< end >>
