magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -1857 244 1857 284
rect -1857 192 -1818 244
rect -1766 192 -1607 244
rect -1555 192 -1397 244
rect -1345 192 -1186 244
rect -1134 192 -975 244
rect -923 192 -764 244
rect -712 192 -553 244
rect -501 192 -343 244
rect -291 192 -132 244
rect -80 192 80 244
rect 132 192 291 244
rect 343 192 501 244
rect 553 192 712 244
rect 764 192 923 244
rect 975 192 1134 244
rect 1186 192 1345 244
rect 1397 192 1555 244
rect 1607 192 1766 244
rect 1818 192 1857 244
rect -1857 26 1857 192
rect -1857 -26 -1818 26
rect -1766 -26 -1607 26
rect -1555 -26 -1397 26
rect -1345 -26 -1186 26
rect -1134 -26 -975 26
rect -923 -26 -764 26
rect -712 -26 -553 26
rect -501 -26 -343 26
rect -291 -26 -132 26
rect -80 -26 80 26
rect 132 -26 291 26
rect 343 -26 501 26
rect 553 -26 712 26
rect 764 -26 923 26
rect 975 -26 1134 26
rect 1186 -26 1345 26
rect 1397 -26 1555 26
rect 1607 -26 1766 26
rect 1818 -26 1857 26
rect -1857 -192 1857 -26
rect -1857 -244 -1818 -192
rect -1766 -244 -1607 -192
rect -1555 -244 -1397 -192
rect -1345 -244 -1186 -192
rect -1134 -244 -975 -192
rect -923 -244 -764 -192
rect -712 -244 -553 -192
rect -501 -244 -343 -192
rect -291 -244 -132 -192
rect -80 -244 80 -192
rect 132 -244 291 -192
rect 343 -244 501 -192
rect 553 -244 712 -192
rect 764 -244 923 -192
rect 975 -244 1134 -192
rect 1186 -244 1345 -192
rect 1397 -244 1555 -192
rect 1607 -244 1766 -192
rect 1818 -244 1857 -192
rect -1857 -284 1857 -244
<< via1 >>
rect -1818 192 -1766 244
rect -1607 192 -1555 244
rect -1397 192 -1345 244
rect -1186 192 -1134 244
rect -975 192 -923 244
rect -764 192 -712 244
rect -553 192 -501 244
rect -343 192 -291 244
rect -132 192 -80 244
rect 80 192 132 244
rect 291 192 343 244
rect 501 192 553 244
rect 712 192 764 244
rect 923 192 975 244
rect 1134 192 1186 244
rect 1345 192 1397 244
rect 1555 192 1607 244
rect 1766 192 1818 244
rect -1818 -26 -1766 26
rect -1607 -26 -1555 26
rect -1397 -26 -1345 26
rect -1186 -26 -1134 26
rect -975 -26 -923 26
rect -764 -26 -712 26
rect -553 -26 -501 26
rect -343 -26 -291 26
rect -132 -26 -80 26
rect 80 -26 132 26
rect 291 -26 343 26
rect 501 -26 553 26
rect 712 -26 764 26
rect 923 -26 975 26
rect 1134 -26 1186 26
rect 1345 -26 1397 26
rect 1555 -26 1607 26
rect 1766 -26 1818 26
rect -1818 -244 -1766 -192
rect -1607 -244 -1555 -192
rect -1397 -244 -1345 -192
rect -1186 -244 -1134 -192
rect -975 -244 -923 -192
rect -764 -244 -712 -192
rect -553 -244 -501 -192
rect -343 -244 -291 -192
rect -132 -244 -80 -192
rect 80 -244 132 -192
rect 291 -244 343 -192
rect 501 -244 553 -192
rect 712 -244 764 -192
rect 923 -244 975 -192
rect 1134 -244 1186 -192
rect 1345 -244 1397 -192
rect 1555 -244 1607 -192
rect 1766 -244 1818 -192
<< metal2 >>
rect -1857 244 1856 284
rect -1857 192 -1818 244
rect -1766 192 -1607 244
rect -1555 192 -1397 244
rect -1345 192 -1186 244
rect -1134 192 -975 244
rect -923 192 -764 244
rect -712 192 -553 244
rect -501 192 -343 244
rect -291 192 -132 244
rect -80 192 80 244
rect 132 192 291 244
rect 343 192 501 244
rect 553 192 712 244
rect 764 192 923 244
rect 975 192 1134 244
rect 1186 192 1345 244
rect 1397 192 1555 244
rect 1607 192 1766 244
rect 1818 192 1856 244
rect -1857 26 1856 192
rect -1857 -26 -1818 26
rect -1766 -26 -1607 26
rect -1555 -26 -1397 26
rect -1345 -26 -1186 26
rect -1134 -26 -975 26
rect -923 -26 -764 26
rect -712 -26 -553 26
rect -501 -26 -343 26
rect -291 -26 -132 26
rect -80 -26 80 26
rect 132 -26 291 26
rect 343 -26 501 26
rect 553 -26 712 26
rect 764 -26 923 26
rect 975 -26 1134 26
rect 1186 -26 1345 26
rect 1397 -26 1555 26
rect 1607 -26 1766 26
rect 1818 -26 1856 26
rect -1857 -192 1856 -26
rect -1857 -244 -1818 -192
rect -1766 -244 -1607 -192
rect -1555 -244 -1397 -192
rect -1345 -244 -1186 -192
rect -1134 -244 -975 -192
rect -923 -244 -764 -192
rect -712 -244 -553 -192
rect -501 -244 -343 -192
rect -291 -244 -132 -192
rect -80 -244 80 -192
rect 132 -244 291 -192
rect 343 -244 501 -192
rect 553 -244 712 -192
rect 764 -244 923 -192
rect 975 -244 1134 -192
rect 1186 -244 1345 -192
rect 1397 -244 1555 -192
rect 1607 -244 1766 -192
rect 1818 -244 1856 -192
rect -1857 -284 1856 -244
<< properties >>
string GDS_END 1063288
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 1059700
<< end >>
