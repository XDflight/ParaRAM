magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -50 230 50 236
rect -50 204 -44 230
rect -18 204 18 230
rect 44 204 50 230
rect -50 168 50 204
rect -50 142 -44 168
rect -18 142 18 168
rect 44 142 50 168
rect -50 106 50 142
rect -50 80 -44 106
rect -18 80 18 106
rect 44 80 50 106
rect -50 44 50 80
rect -50 18 -44 44
rect -18 18 18 44
rect 44 18 50 44
rect -50 -18 50 18
rect -50 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 50 -18
rect -50 -80 50 -44
rect -50 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 50 -80
rect -50 -142 50 -106
rect -50 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 50 -142
rect -50 -204 50 -168
rect -50 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 50 -204
rect -50 -236 50 -230
<< via1 >>
rect -44 204 -18 230
rect 18 204 44 230
rect -44 142 -18 168
rect 18 142 44 168
rect -44 80 -18 106
rect 18 80 44 106
rect -44 18 -18 44
rect 18 18 44 44
rect -44 -44 -18 -18
rect 18 -44 44 -18
rect -44 -106 -18 -80
rect 18 -106 44 -80
rect -44 -168 -18 -142
rect 18 -168 44 -142
rect -44 -230 -18 -204
rect 18 -230 44 -204
<< metal2 >>
rect -50 230 50 236
rect -50 204 -44 230
rect -18 204 18 230
rect 44 204 50 230
rect -50 168 50 204
rect -50 142 -44 168
rect -18 142 18 168
rect 44 142 50 168
rect -50 106 50 142
rect -50 80 -44 106
rect -18 80 18 106
rect 44 80 50 106
rect -50 44 50 80
rect -50 18 -44 44
rect -18 18 18 44
rect 44 18 50 44
rect -50 -18 50 18
rect -50 -44 -44 -18
rect -18 -44 18 -18
rect 44 -44 50 -18
rect -50 -80 50 -44
rect -50 -106 -44 -80
rect -18 -106 18 -80
rect 44 -106 50 -80
rect -50 -142 50 -106
rect -50 -168 -44 -142
rect -18 -168 18 -142
rect 44 -168 50 -142
rect -50 -204 50 -168
rect -50 -230 -44 -204
rect -18 -230 18 -204
rect 44 -230 50 -204
rect -50 -236 50 -230
<< properties >>
string GDS_END 526944
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 525788
<< end >>
