magic
tech gf180mcuB
magscale 1 5
timestamp 1666464484
<< metal3 >>
rect 357 911 857 1215
use M2_M143105899832101_64x8m81  M2_M143105899832101_64x8m81_0
timestamp 1666464484
transform 1 0 607 0 1 993
box -236 -81 236 81
use M3_M243105899832100_64x8m81  M3_M243105899832100_64x8m81_0
timestamp 1666464484
transform 1 0 607 0 1 993
box -236 -81 236 81
<< properties >>
string GDS_END 2272246
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 2272074
<< end >>
