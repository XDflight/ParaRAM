magic
tech gf180mcuC
magscale 1 5
timestamp 1666464484
<< metal1 >>
rect -143 44 143 50
rect -143 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 143 44
rect -143 -18 143 18
rect -143 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 143 -18
rect -143 -50 143 -44
<< via1 >>
rect -137 18 -111 44
rect -75 18 -49 44
rect -13 18 13 44
rect 49 18 75 44
rect 111 18 137 44
rect -137 -44 -111 -18
rect -75 -44 -49 -18
rect -13 -44 13 -18
rect 49 -44 75 -18
rect 111 -44 137 -18
<< metal2 >>
rect -143 44 143 50
rect -143 18 -137 44
rect -111 18 -75 44
rect -49 18 -13 44
rect 13 18 49 44
rect 75 18 111 44
rect 137 18 143 44
rect -143 -18 143 18
rect -143 -44 -137 -18
rect -111 -44 -75 -18
rect -49 -44 -13 -18
rect 13 -44 49 -18
rect 75 -44 111 -18
rect 137 -44 143 -18
rect -143 -50 143 -44
<< properties >>
string GDS_END 2145014
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 2144242
<< end >>
