magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -203 10266 787 12370
rect -7 8752 622 10266
rect -7 8695 624 8752
rect -5 7108 624 8695
rect -5 1620 624 3202
rect -221 1164 756 1620
rect -203 648 756 1164
<< pmos >>
rect 138 11191 258 11873
rect 362 11191 482 11873
rect 138 10416 258 11098
rect 362 10416 482 11098
rect 67 788 187 1085
rect 319 788 439 1085
<< pdiff >>
rect -67 11828 138 11873
rect -67 11782 -23 11828
rect 23 11782 138 11828
rect -67 11646 138 11782
rect -67 11600 -23 11646
rect 23 11600 138 11646
rect -67 11465 138 11600
rect -67 11419 -23 11465
rect 23 11419 138 11465
rect -67 11283 138 11419
rect -67 11237 -23 11283
rect 23 11237 138 11283
rect -67 11191 138 11237
rect 258 11828 362 11873
rect 258 11782 287 11828
rect 333 11782 362 11828
rect 258 11646 362 11782
rect 258 11600 287 11646
rect 333 11600 362 11646
rect 258 11465 362 11600
rect 258 11419 287 11465
rect 333 11419 362 11465
rect 258 11283 362 11419
rect 258 11237 287 11283
rect 333 11237 362 11283
rect 258 11191 362 11237
rect 482 11828 650 11873
rect 482 11782 513 11828
rect 559 11782 650 11828
rect 482 11646 650 11782
rect 482 11600 513 11646
rect 559 11600 650 11646
rect 482 11465 650 11600
rect 482 11419 513 11465
rect 559 11419 650 11465
rect 482 11283 650 11419
rect 482 11237 513 11283
rect 559 11237 650 11283
rect 482 11191 650 11237
rect -67 11052 138 11098
rect -67 11006 -23 11052
rect 23 11006 138 11052
rect -67 10871 138 11006
rect -67 10825 -23 10871
rect 23 10825 138 10871
rect -67 10690 138 10825
rect -67 10644 -23 10690
rect 23 10644 138 10690
rect -67 10508 138 10644
rect -67 10462 -23 10508
rect 23 10462 138 10508
rect -67 10416 138 10462
rect 258 11052 362 11098
rect 258 11006 287 11052
rect 333 11006 362 11052
rect 258 10871 362 11006
rect 258 10825 287 10871
rect 333 10825 362 10871
rect 258 10690 362 10825
rect 258 10644 287 10690
rect 333 10644 362 10690
rect 258 10508 362 10644
rect 258 10462 287 10508
rect 333 10462 362 10508
rect 258 10416 362 10462
rect 482 11052 650 11098
rect 482 11006 513 11052
rect 559 11006 650 11052
rect 482 10871 650 11006
rect 482 10825 513 10871
rect 559 10825 650 10871
rect 482 10690 650 10825
rect 482 10644 513 10690
rect 559 10644 650 10690
rect 482 10508 650 10644
rect 482 10462 513 10508
rect 559 10462 650 10508
rect 482 10416 650 10462
rect -67 960 67 1085
rect -67 914 -23 960
rect 23 914 67 960
rect -67 788 67 914
rect 187 960 319 1085
rect 187 914 230 960
rect 276 914 319 960
rect 187 788 319 914
rect 439 960 620 1085
rect 439 914 480 960
rect 526 914 620 960
rect 439 788 620 914
<< pdiffc >>
rect -23 11782 23 11828
rect -23 11600 23 11646
rect -23 11419 23 11465
rect -23 11237 23 11283
rect 287 11782 333 11828
rect 287 11600 333 11646
rect 287 11419 333 11465
rect 287 11237 333 11283
rect 513 11782 559 11828
rect 513 11600 559 11646
rect 513 11419 559 11465
rect 513 11237 559 11283
rect -23 11006 23 11052
rect -23 10825 23 10871
rect -23 10644 23 10690
rect -23 10462 23 10508
rect 287 11006 333 11052
rect 287 10825 333 10871
rect 287 10644 333 10690
rect 287 10462 333 10508
rect 513 11006 559 11052
rect 513 10825 559 10871
rect 513 10644 559 10690
rect 513 10462 559 10508
rect -23 914 23 960
rect 230 914 276 960
rect 480 914 526 960
<< psubdiff >>
rect -80 5260 80 5320
rect -80 5214 -23 5260
rect 23 5214 80 5260
rect -80 5154 80 5214
rect 14 164 474 183
rect 14 118 33 164
rect 455 118 474 164
rect 14 99 474 118
<< nsubdiff >>
rect -1 12165 650 12222
rect -1 12119 129 12165
rect 175 12119 287 12165
rect 333 12119 445 12165
rect 491 12119 650 12165
rect -1 12062 650 12119
rect -78 1415 620 1472
rect -78 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -78 1312 620 1369
<< psubdiffcont >>
rect -23 5214 23 5260
rect 33 118 455 164
<< nsubdiffcont >>
rect 129 12119 175 12165
rect 287 12119 333 12165
rect 445 12119 491 12165
rect -23 1369 23 1415
rect 135 1369 181 1415
rect 293 1369 339 1415
rect 451 1369 497 1415
<< polysilicon >>
rect 138 11873 258 11946
rect 362 11873 482 11946
rect 138 11098 258 11191
rect 362 11098 482 11191
rect 138 10356 258 10416
rect 362 10356 482 10416
rect 138 10334 482 10356
rect 138 10288 234 10334
rect 374 10288 482 10334
rect 138 10269 482 10288
rect 248 10198 368 10269
rect 250 7167 370 7249
rect 250 7121 287 7167
rect 333 7121 370 7167
rect 250 7102 370 7121
rect 250 4887 370 5558
rect 250 3469 370 3554
rect 250 3423 287 3469
rect 333 3423 370 3469
rect 250 3404 370 3423
rect 250 3192 370 3211
rect 250 3146 287 3192
rect 333 3146 370 3192
rect 250 3061 370 3146
rect 67 1225 439 1244
rect 67 1179 230 1225
rect 276 1179 439 1225
rect 67 1145 439 1179
rect 67 1085 187 1145
rect 319 1085 439 1145
rect 67 619 187 788
rect 67 612 186 619
rect 66 539 186 612
rect 319 601 439 788
rect 319 570 410 601
rect 290 539 410 570
rect 66 497 184 498
rect 66 310 186 382
rect 290 310 410 382
<< polycontact >>
rect 234 10288 374 10334
rect 287 7121 333 7167
rect 287 3423 333 3469
rect 287 3146 333 3192
rect 230 1179 276 1225
<< metal1 >>
rect -58 12203 620 12227
rect -58 12165 281 12203
rect 333 12165 620 12203
rect -58 12119 129 12165
rect 175 12151 281 12165
rect 175 12119 287 12151
rect 333 12119 445 12165
rect 491 12119 620 12165
rect -58 12017 620 12119
rect -58 11965 281 12017
rect 333 11965 620 12017
rect -58 11944 620 11965
rect -58 11828 147 11944
rect -58 11782 -23 11828
rect 23 11782 147 11828
rect -58 11646 147 11782
rect -58 11600 -23 11646
rect 23 11600 147 11646
rect -58 11465 147 11600
rect -58 11419 -23 11465
rect 23 11419 147 11465
rect -58 11283 147 11419
rect -58 11237 -23 11283
rect 23 11237 147 11283
rect -58 11052 147 11237
rect 252 11828 367 11864
rect 252 11782 287 11828
rect 333 11782 367 11828
rect 252 11646 367 11782
rect 252 11613 287 11646
rect 252 11457 264 11613
rect 333 11600 367 11646
rect 316 11465 367 11600
rect 252 11419 287 11457
rect 333 11419 367 11465
rect 252 11283 367 11419
rect 252 11237 287 11283
rect 333 11237 367 11283
rect 252 11200 367 11237
rect 472 11828 620 11944
rect 472 11782 513 11828
rect 559 11782 620 11828
rect 472 11646 620 11782
rect 472 11600 513 11646
rect 559 11600 620 11646
rect 472 11465 620 11600
rect 472 11419 513 11465
rect 559 11419 620 11465
rect 472 11283 620 11419
rect 472 11237 513 11283
rect 559 11237 620 11283
rect -58 11006 -23 11052
rect 23 11006 147 11052
rect -58 10871 147 11006
rect -58 10825 -23 10871
rect 23 10825 147 10871
rect -58 10690 147 10825
rect -58 10644 -23 10690
rect 23 10644 147 10690
rect -58 10508 147 10644
rect -58 10462 -23 10508
rect 23 10462 147 10508
rect -58 10425 147 10462
rect 252 11052 367 11089
rect 252 11006 287 11052
rect 333 11006 367 11052
rect 252 10871 367 11006
rect 252 10825 287 10871
rect 333 10834 367 10871
rect 252 10690 303 10825
rect 252 10644 287 10690
rect 355 10678 367 10834
rect 333 10644 367 10678
rect 252 10508 367 10644
rect 252 10462 287 10508
rect 333 10462 367 10508
rect 252 10425 367 10462
rect 472 11052 620 11237
rect 472 11006 513 11052
rect 559 11006 620 11052
rect 472 10871 620 11006
rect 472 10825 513 10871
rect 559 10825 620 10871
rect 472 10690 620 10825
rect 472 10644 513 10690
rect 559 10644 620 10690
rect 472 10508 620 10644
rect 472 10462 513 10508
rect 559 10462 620 10508
rect 472 10425 620 10462
rect 78 10334 453 10345
rect 78 10288 234 10334
rect 374 10288 453 10334
rect 78 10271 453 10288
rect 58 9646 219 9658
rect 58 9490 70 9646
rect 122 9490 219 9646
rect 58 9478 219 9490
rect 397 9646 558 9658
rect 397 9490 494 9646
rect 546 9490 558 9646
rect 397 9478 558 9490
rect 67 8598 177 8610
rect 67 8442 79 8598
rect 131 8442 177 8598
rect 67 8430 177 8442
rect 70 7248 177 8430
rect 433 7248 549 8610
rect 70 6919 141 7248
rect 219 7167 400 7178
rect 219 7121 287 7167
rect 333 7163 400 7167
rect 219 7007 301 7121
rect 353 7007 400 7163
rect 219 6995 400 7007
rect 479 6919 549 7248
rect 70 5557 184 6919
rect 443 5657 549 6919
rect 364 5567 549 5657
rect 364 5487 457 5567
rect 45 5483 457 5487
rect -154 5463 457 5483
rect -154 5411 -114 5463
rect -62 5411 72 5463
rect 124 5411 457 5463
rect -154 5391 457 5411
rect 45 5390 457 5391
rect -71 5306 71 5311
rect -71 5265 620 5306
rect -71 5260 114 5265
rect -71 5214 -23 5260
rect 23 5214 114 5260
rect -71 5213 114 5214
rect 166 5213 620 5265
rect -71 5172 620 5213
rect -71 5163 71 5172
rect 48 5061 561 5084
rect 48 5009 494 5061
rect 546 5009 561 5061
rect 48 4987 561 5009
rect 48 4915 141 4987
rect 48 3568 188 4915
rect 48 3553 192 3568
rect 443 3553 549 4915
rect 48 3060 141 3553
rect 219 3469 400 3483
rect 219 3423 287 3469
rect 333 3423 400 3469
rect 219 3420 400 3423
rect 219 3368 286 3420
rect 338 3368 400 3420
rect 219 3348 400 3368
rect 219 3225 400 3268
rect 219 3173 232 3225
rect 388 3173 400 3225
rect 219 3146 287 3173
rect 333 3146 400 3173
rect 219 3132 400 3146
rect 479 3060 549 3553
rect 48 1708 181 3060
rect 435 1710 549 3060
rect 364 1554 549 1710
rect -58 1415 620 1452
rect -58 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -58 1332 620 1369
rect -57 960 57 1332
rect 136 1229 445 1252
rect 136 1225 355 1229
rect 136 1179 230 1225
rect 276 1179 355 1225
rect 136 1177 355 1179
rect 407 1177 445 1229
rect 136 1155 445 1177
rect 549 1076 620 1332
rect -57 914 -23 960
rect 23 914 57 960
rect -57 797 57 914
rect 195 1064 323 1076
rect 195 908 207 1064
rect 259 960 323 1064
rect 276 914 323 960
rect 259 908 323 914
rect 195 797 323 908
rect 446 960 620 1076
rect 446 914 480 960
rect 526 914 620 960
rect 446 797 620 914
rect -58 271 57 500
rect 215 380 288 797
rect 439 271 620 500
rect -58 164 620 271
rect -58 118 33 164
rect 455 118 620 164
rect -58 76 620 118
<< via1 >>
rect 281 12165 333 12203
rect 281 12151 287 12165
rect 287 12151 333 12165
rect 281 11965 333 12017
rect 264 11600 287 11613
rect 287 11600 316 11613
rect 264 11465 316 11600
rect 264 11457 287 11465
rect 287 11457 316 11465
rect 303 10825 333 10834
rect 333 10825 355 10834
rect 303 10690 355 10825
rect 303 10678 333 10690
rect 333 10678 355 10690
rect 70 9490 122 9646
rect 494 9490 546 9646
rect 79 8442 131 8598
rect 301 7121 333 7163
rect 333 7121 353 7163
rect 301 7007 353 7121
rect -114 5411 -62 5463
rect 72 5411 124 5463
rect 114 5213 166 5265
rect 494 5009 546 5061
rect 286 3368 338 3420
rect 232 3192 388 3225
rect 232 3173 287 3192
rect 287 3173 333 3192
rect 333 3173 388 3192
rect 355 1177 407 1229
rect 207 960 259 1064
rect 207 914 230 960
rect 230 914 259 960
rect 207 908 259 914
<< metal2 >>
rect 77 11563 133 12370
rect 246 12205 374 12227
rect 246 12149 279 12205
rect 335 12149 374 12205
rect 246 12019 374 12149
rect 246 11963 279 12019
rect 335 11963 374 12019
rect 246 11944 374 11963
rect 252 11613 328 11625
rect 252 11563 264 11613
rect 77 11507 264 11563
rect 77 9658 133 11507
rect 252 11457 264 11507
rect 316 11457 328 11613
rect 252 11445 328 11457
rect 291 10834 367 10846
rect 291 10678 303 10834
rect 355 10784 367 10834
rect 492 10784 548 12370
rect 355 10728 548 10784
rect 355 10678 367 10728
rect 291 10666 367 10678
rect 492 9658 548 10728
rect 58 9646 134 9658
rect 58 9490 70 9646
rect 122 9490 134 9646
rect 58 9478 134 9490
rect 482 9646 558 9658
rect 482 9490 494 9646
rect 546 9490 558 9646
rect 482 9478 558 9490
rect 77 8610 133 9478
rect 67 8598 143 8610
rect 67 8442 79 8598
rect 131 8442 143 8598
rect 67 8430 143 8442
rect 77 5585 133 8430
rect 289 7163 365 7175
rect 289 7007 301 7163
rect 353 7007 365 7163
rect 289 6995 365 7007
rect -154 5463 154 5483
rect -154 5411 -114 5463
rect -62 5411 72 5463
rect 124 5411 154 5463
rect -154 5391 154 5411
rect -154 -1 -66 5391
rect 76 5267 205 5306
rect 76 5211 112 5267
rect 168 5211 205 5267
rect 76 5172 205 5211
rect 76 5049 204 5172
rect 76 4993 112 5049
rect 168 4993 204 5049
rect 76 4955 204 4993
rect 299 4812 355 6995
rect 492 5073 548 9478
rect 482 5061 558 5073
rect 482 5009 494 5061
rect 546 5009 558 5061
rect 482 4997 558 5009
rect 81 4756 355 4812
rect 81 3237 137 4756
rect 250 3420 573 3444
rect 250 3368 286 3420
rect 338 3368 573 3420
rect 250 3347 573 3368
rect 81 3225 400 3237
rect 81 3173 232 3225
rect 388 3173 400 3225
rect 81 3161 400 3173
rect 81 1076 137 3161
rect 481 1853 573 3347
rect 382 1756 573 1853
rect 382 1252 475 1756
rect 316 1229 475 1252
rect 316 1177 355 1229
rect 407 1177 475 1229
rect 316 1155 475 1177
rect 81 1064 271 1076
rect 81 1020 207 1064
rect 195 908 207 1020
rect 259 908 271 1064
rect 195 896 271 908
rect 246 49 374 278
<< via2 >>
rect 279 12203 335 12205
rect 279 12151 281 12203
rect 281 12151 333 12203
rect 333 12151 335 12203
rect 279 12149 335 12151
rect 279 12017 335 12019
rect 279 11965 281 12017
rect 281 11965 333 12017
rect 333 11965 335 12017
rect 279 11963 335 11965
rect 112 5265 168 5267
rect 112 5213 114 5265
rect 114 5213 166 5265
rect 166 5213 168 5265
rect 112 5211 168 5213
rect 112 4993 168 5049
<< metal3 >>
rect -65 12205 929 12347
rect -65 12149 279 12205
rect 335 12149 929 12205
rect -65 12019 929 12149
rect -65 11963 279 12019
rect 335 11963 929 12019
rect -65 10538 929 11963
rect -1 5267 930 6537
rect -1 5211 112 5267
rect 168 5211 930 5267
rect -1 5049 930 5211
rect -1 4993 112 5049
rect 168 4993 930 5049
rect -1 4657 930 4993
rect -1 4331 929 4546
rect -1 4009 929 4224
rect -1 3688 929 3903
rect -1 3366 929 3581
rect -1 2674 929 2889
rect -1 2352 929 2567
rect -1 2030 929 2245
rect -1 1708 929 1923
rect -1 1160 929 1602
rect -1 49 929 504
use M1_NWELL$$46277676_256x8m81_0  M1_NWELL$$46277676_256x8m81_0_0
timestamp 1666464484
transform 1 0 310 0 1 12142
box 0 0 1 1
use M1_NWELL$$47121452_256x8m81_0  M1_NWELL$$47121452_256x8m81_0_0
timestamp 1666464484
transform 1 0 237 0 1 1392
box 0 0 1 1
use M1_PACTIVE4310590878140_256x8m81  M1_PACTIVE4310590878140_256x8m81_0
timestamp 1666464484
transform 1 0 244 0 1 141
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_0
timestamp 1666464484
transform 1 0 310 0 1 3446
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_1
timestamp 1666464484
transform 1 0 310 0 1 3169
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_2
timestamp 1666464484
transform 1 0 253 0 1 1202
box 0 0 1 1
use M1_POLY24310590878127_256x8m81  M1_POLY24310590878127_256x8m81_3
timestamp 1666464484
transform 1 0 310 0 1 7144
box 0 0 1 1
use M1_POLY24310590878129_256x8m81  M1_POLY24310590878129_256x8m81_0
timestamp 1666464484
transform 1 0 304 0 1 10311
box 0 0 1 1
use M1_PSUB$$45111340_256x8m81_0  M1_PSUB$$45111340_256x8m81_0_0
timestamp 1666464484
transform 1 0 0 0 1 5237
box 0 0 1 1
use M2_M1$$46894124_256x8m81_0  M2_M1$$46894124_256x8m81_0_0
timestamp 1666464484
transform 1 0 140 0 1 5239
box 0 0 1 1
use M2_M14310590878116_256x8m81  M2_M14310590878116_256x8m81_0
timestamp 1666464484
transform 1 0 520 0 1 5035
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_0
timestamp 1666464484
transform 0 1 310 -1 0 3199
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_1
timestamp 1666464484
transform 1 0 96 0 1 9568
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_2
timestamp 1666464484
transform 1 0 329 0 1 10756
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_3
timestamp 1666464484
transform 1 0 290 0 1 11535
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_4
timestamp 1666464484
transform 1 0 105 0 1 8520
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_5
timestamp 1666464484
transform 1 0 233 0 1 986
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_6
timestamp 1666464484
transform 1 0 327 0 1 7085
box 0 0 1 1
use M2_M14310590878119_256x8m81  M2_M14310590878119_256x8m81_7
timestamp 1666464484
transform 1 0 520 0 1 9568
box 0 0 1 1
use M3_M2$$43368492_256x8m81  M3_M2$$43368492_256x8m81_0
timestamp 1666464484
transform 1 0 140 0 1 5130
box 0 0 1 1
use nmos_5p0431059087811_256x8m81  nmos_5p0431059087811_256x8m81_0
timestamp 1666464484
transform 1 0 66 0 1 383
box -88 -44 432 158
use nmos_5p0431059087812_256x8m81  nmos_5p0431059087812_256x8m81_0
timestamp 1666464484
transform 1 0 250 0 -1 6919
box -88 -44 208 1406
use nmos_5p0431059087812_256x8m81  nmos_5p0431059087812_256x8m81_1
timestamp 1666464484
transform 1 0 250 0 -1 4915
box -88 -44 208 1406
use pmos_5p0431059087810_256x8m81  pmos_5p0431059087810_256x8m81_0
timestamp 1666464484
transform 1 0 250 0 -1 3060
box -208 -120 328 1482
use pmos_5p0431059087810_256x8m81  pmos_5p0431059087810_256x8m81_1
timestamp 1666464484
transform 1 0 248 0 -1 10197
box -208 -120 328 1482
use pmos_5p0431059087810_256x8m81  pmos_5p0431059087810_256x8m81_2
timestamp 1666464484
transform 1 0 250 0 -1 8610
box -208 -120 328 1482
use via1_2_256x8m81_0  via1_2_256x8m81_0_0
timestamp 1666464484
transform 1 0 264 0 1 88
box -1 -1 93 128
use via1_R90_256x8m81_0  via1_R90_256x8m81_0_0
timestamp 1666464484
transform 0 -1 378 1 0 3348
box 0 0 1 1
use via1_R90_256x8m81_0  via1_R90_256x8m81_0_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
use via1_R90_256x8m81_0  via1_R90_256x8m81_0_2
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via1_R270_256x8m81_0  via1_R270_256x8m81_0_0
timestamp 1666464484
transform 0 1 317 -1 0 1251
box 0 0 1 1
use via1_x2_R90_256x8m81_0  via1_x2_R90_256x8m81_0_0
timestamp 1666464484
transform 0 1 -154 1 0 5391
box 0 0 1 1
use via2_R90_256x8m81_0  via2_R90_256x8m81_0_0
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_256x8m81_0  via2_R90_256x8m81_0_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
<< labels >>
rlabel metal1 s 492 1805 492 1805 4 d
port 1 nsew
rlabel metal1 s 259 10272 259 10272 4 pcb
port 2 nsew
rlabel metal1 s 318 1356 318 1356 4 vdd
port 3 nsew
rlabel metal3 s 279 91 279 91 4 vss
port 4 nsew
rlabel metal3 s 318 12094 318 12094 4 vdd
port 3 nsew
rlabel metal3 s 303 5255 303 5255 4 vss
port 4 nsew
rlabel metal2 s 518 11931 518 11931 4 b
port 5 nsew
rlabel metal2 s 105 11931 105 11931 4 bb
port 6 nsew
rlabel metal2 s 0 304 0 304 4 db
port 7 nsew
rlabel metal2 s 285 1222 285 1222 4 ypass
port 8 nsew
<< properties >>
string GDS_END 515262
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 505852
string path 0.525 61.850 0.525 27.925 
<< end >>
