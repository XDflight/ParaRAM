magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect -170 1005 170 1046
rect -170 953 -132 1005
rect -80 953 80 1005
rect 132 953 170 1005
rect -170 788 170 953
rect -170 736 -132 788
rect -80 736 80 788
rect 132 736 170 788
rect -170 570 170 736
rect -170 518 -132 570
rect -80 518 80 570
rect 132 518 170 570
rect -170 353 170 518
rect -170 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -170 135 170 301
rect -170 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -170 -83 170 83
rect -170 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -170 -301 170 -135
rect -170 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -170 -518 170 -353
rect -170 -570 -132 -518
rect -80 -570 80 -518
rect 132 -570 170 -518
rect -170 -736 170 -570
rect -170 -788 -132 -736
rect -80 -788 80 -736
rect 132 -788 170 -736
rect -170 -953 170 -788
rect -170 -1005 -132 -953
rect -80 -1005 80 -953
rect 132 -1005 170 -953
rect -170 -1046 170 -1005
<< via1 >>
rect -132 953 -80 1005
rect 80 953 132 1005
rect -132 736 -80 788
rect 80 736 132 788
rect -132 518 -80 570
rect 80 518 132 570
rect -132 301 -80 353
rect 80 301 132 353
rect -132 83 -80 135
rect 80 83 132 135
rect -132 -135 -80 -83
rect 80 -135 132 -83
rect -132 -353 -80 -301
rect 80 -353 132 -301
rect -132 -570 -80 -518
rect 80 -570 132 -518
rect -132 -788 -80 -736
rect 80 -788 132 -736
rect -132 -1005 -80 -953
rect 80 -1005 132 -953
<< metal2 >>
rect -170 1005 170 1046
rect -170 953 -132 1005
rect -80 953 80 1005
rect 132 953 170 1005
rect -170 788 170 953
rect -170 736 -132 788
rect -80 736 80 788
rect 132 736 170 788
rect -170 570 170 736
rect -170 518 -132 570
rect -80 518 80 570
rect 132 518 170 570
rect -170 353 170 518
rect -170 301 -132 353
rect -80 301 80 353
rect 132 301 170 353
rect -170 135 170 301
rect -170 83 -132 135
rect -80 83 80 135
rect 132 83 170 135
rect -170 -83 170 83
rect -170 -135 -132 -83
rect -80 -135 80 -83
rect 132 -135 170 -83
rect -170 -301 170 -135
rect -170 -353 -132 -301
rect -80 -353 80 -301
rect 132 -353 170 -301
rect -170 -518 170 -353
rect -170 -570 -132 -518
rect -80 -570 80 -518
rect 132 -570 170 -518
rect -170 -736 170 -570
rect -170 -788 -132 -736
rect -80 -788 80 -736
rect 132 -788 170 -736
rect -170 -953 170 -788
rect -170 -1005 -132 -953
rect -80 -1005 80 -953
rect 132 -1005 170 -953
rect -170 -1046 170 -1005
<< properties >>
string GDS_END 896960
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 895548
<< end >>
