magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< psubdiff >>
rect -1108 23 1108 83
rect -1108 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1108 23
rect -1108 -83 1108 -23
<< psubdiffcont >>
rect -1051 -23 -1005 23
rect -893 -23 -847 23
rect -735 -23 -689 23
rect -577 -23 -531 23
rect -418 -23 -372 23
rect -260 -23 -214 23
rect -102 -23 -56 23
rect 56 -23 102 23
rect 214 -23 260 23
rect 372 -23 418 23
rect 531 -23 577 23
rect 689 -23 735 23
rect 847 -23 893 23
rect 1005 -23 1051 23
<< metal1 >>
rect -1099 23 1099 74
rect -1099 -23 -1051 23
rect -1005 -23 -893 23
rect -847 -23 -735 23
rect -689 -23 -577 23
rect -531 -23 -418 23
rect -372 -23 -260 23
rect -214 -23 -102 23
rect -56 -23 56 23
rect 102 -23 214 23
rect 260 -23 372 23
rect 418 -23 531 23
rect 577 -23 689 23
rect 735 -23 847 23
rect 893 -23 1005 23
rect 1051 -23 1099 23
rect -1099 -74 1099 -23
<< properties >>
string GDS_END 337110
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 336018
<< end >>
