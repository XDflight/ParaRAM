magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -286 -141 344 1275
<< polysilicon >>
rect -31 1135 89 1196
rect -30 -74 88 -1
use pmos_5p04310590548765_128x8m81  pmos_5p04310590548765_128x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -208 -120 328 1274
<< properties >>
string GDS_END 367058
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 366744
<< end >>
