magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 377 5126 870
rect -86 352 1291 377
rect 1975 352 2594 377
rect 3730 352 5126 377
<< pwell >>
rect 1291 352 1975 377
rect 2594 352 3730 377
rect -86 -86 5126 352
<< mvnmos >>
rect 124 156 244 228
rect 348 156 468 228
rect 516 156 636 228
rect 740 156 860 228
rect 908 156 1028 228
rect 1185 135 1305 228
rect 1648 139 1768 232
rect 2060 124 2180 196
rect 2284 124 2404 196
rect 2488 124 2608 196
rect 2788 185 2908 257
rect 2956 185 3076 257
rect 3180 185 3300 257
rect 3404 185 3524 257
rect 3885 106 4005 178
rect 4110 106 4230 178
rect 4370 106 4490 199
rect 4738 68 4858 232
<< mvpmos >>
rect 124 502 224 628
rect 348 502 448 628
rect 496 502 596 628
rect 740 502 840 628
rect 888 502 988 628
rect 1185 502 1285 687
rect 1648 497 1748 660
rect 1996 497 2096 622
rect 2236 474 2336 599
rect 2476 516 2576 641
rect 2768 516 2868 641
rect 2976 516 3076 641
rect 3377 503 3477 628
rect 3581 503 3681 628
rect 3982 527 4082 652
rect 4186 527 4286 652
rect 4426 527 4526 712
rect 4778 472 4878 716
<< mvndiff >>
rect 1365 244 1437 257
rect 1365 228 1378 244
rect 36 215 124 228
rect 36 169 49 215
rect 95 169 124 215
rect 36 156 124 169
rect 244 215 348 228
rect 244 169 273 215
rect 319 169 348 215
rect 244 156 348 169
rect 468 156 516 228
rect 636 215 740 228
rect 636 169 665 215
rect 711 169 740 215
rect 636 156 740 169
rect 860 156 908 228
rect 1028 194 1185 228
rect 1028 156 1110 194
rect 1097 148 1110 156
rect 1156 148 1185 194
rect 1097 135 1185 148
rect 1305 198 1378 228
rect 1424 198 1437 244
rect 1828 244 1900 257
rect 1828 232 1841 244
rect 1305 135 1437 198
rect 1560 198 1648 232
rect 1560 152 1573 198
rect 1619 152 1648 198
rect 1560 139 1648 152
rect 1768 198 1841 232
rect 1887 198 1900 244
rect 1768 139 1900 198
rect 2668 196 2788 257
rect 1972 183 2060 196
rect 1972 137 1985 183
rect 2031 137 2060 183
rect 1972 124 2060 137
rect 2180 183 2284 196
rect 2180 137 2209 183
rect 2255 137 2284 183
rect 2180 124 2284 137
rect 2404 124 2488 196
rect 2608 185 2788 196
rect 2908 185 2956 257
rect 3076 244 3180 257
rect 3076 198 3105 244
rect 3151 198 3180 244
rect 3076 185 3180 198
rect 3300 244 3404 257
rect 3300 198 3329 244
rect 3375 198 3404 244
rect 3300 185 3404 198
rect 3524 244 3612 257
rect 3524 198 3553 244
rect 3599 198 3612 244
rect 3524 185 3612 198
rect 2608 183 2728 185
rect 2608 137 2637 183
rect 2683 137 2728 183
rect 4290 178 4370 199
rect 3797 165 3885 178
rect 2608 124 2728 137
rect 3797 119 3810 165
rect 3856 119 3885 165
rect 3797 106 3885 119
rect 4005 106 4110 178
rect 4230 165 4370 178
rect 4230 119 4295 165
rect 4341 119 4370 165
rect 4230 106 4370 119
rect 4490 186 4578 199
rect 4490 140 4519 186
rect 4565 140 4578 186
rect 4490 106 4578 140
rect 4650 142 4738 232
rect 4650 96 4663 142
rect 4709 96 4738 142
rect 4650 68 4738 96
rect 4858 177 4946 232
rect 4858 131 4887 177
rect 4933 131 4946 177
rect 4858 68 4946 131
<< mvpdiff >>
rect 1516 716 1588 729
rect 1048 634 1185 687
rect 1048 628 1075 634
rect 36 585 124 628
rect 36 539 49 585
rect 95 539 124 585
rect 36 502 124 539
rect 224 615 348 628
rect 224 569 263 615
rect 309 569 348 615
rect 224 502 348 569
rect 448 502 496 628
rect 596 595 740 628
rect 596 549 665 595
rect 711 549 740 595
rect 596 502 740 549
rect 840 502 888 628
rect 988 588 1075 628
rect 1121 588 1185 634
rect 988 502 1185 588
rect 1285 561 1393 687
rect 1285 515 1322 561
rect 1368 515 1393 561
rect 1285 502 1393 515
rect 1516 670 1529 716
rect 1575 670 1588 716
rect 1516 660 1588 670
rect 2636 735 2708 748
rect 2636 689 2649 735
rect 2695 689 2708 735
rect 1516 497 1648 660
rect 1748 559 1836 660
rect 2636 641 2708 689
rect 1748 513 1777 559
rect 1823 513 1836 559
rect 1748 497 1836 513
rect 1908 571 1996 622
rect 1908 525 1921 571
rect 1967 525 1996 571
rect 1908 497 1996 525
rect 2096 599 2176 622
rect 2396 599 2476 641
rect 2096 562 2236 599
rect 2096 516 2160 562
rect 2206 516 2236 562
rect 2096 497 2236 516
rect 2156 474 2236 497
rect 2336 516 2476 599
rect 2576 516 2768 641
rect 2868 575 2976 641
rect 2868 529 2897 575
rect 2943 529 2976 575
rect 2868 516 2976 529
rect 3076 628 3164 641
rect 4346 652 4426 712
rect 3892 639 3982 652
rect 3076 582 3105 628
rect 3151 582 3164 628
rect 3076 516 3164 582
rect 3289 566 3377 628
rect 3289 520 3302 566
rect 3348 520 3377 566
rect 2336 474 2416 516
rect 3289 503 3377 520
rect 3477 583 3581 628
rect 3477 537 3506 583
rect 3552 537 3581 583
rect 3477 503 3581 537
rect 3681 562 3773 628
rect 3681 516 3710 562
rect 3756 516 3773 562
rect 3892 593 3905 639
rect 3951 593 3982 639
rect 3892 527 3982 593
rect 4082 586 4186 652
rect 4082 540 4111 586
rect 4157 540 4186 586
rect 4082 527 4186 540
rect 4286 639 4426 652
rect 4286 593 4329 639
rect 4375 593 4426 639
rect 4286 527 4426 593
rect 4526 590 4614 712
rect 4526 544 4555 590
rect 4601 544 4614 590
rect 4526 527 4614 544
rect 4690 665 4778 716
rect 3681 503 3773 516
rect 4690 525 4703 665
rect 4749 525 4778 665
rect 4690 472 4778 525
rect 4878 665 4966 716
rect 4878 525 4907 665
rect 4953 525 4966 665
rect 4878 472 4966 525
<< mvndiffc >>
rect 49 169 95 215
rect 273 169 319 215
rect 665 169 711 215
rect 1110 148 1156 194
rect 1378 198 1424 244
rect 1573 152 1619 198
rect 1841 198 1887 244
rect 1985 137 2031 183
rect 2209 137 2255 183
rect 3105 198 3151 244
rect 3329 198 3375 244
rect 3553 198 3599 244
rect 2637 137 2683 183
rect 3810 119 3856 165
rect 4295 119 4341 165
rect 4519 140 4565 186
rect 4663 96 4709 142
rect 4887 131 4933 177
<< mvpdiffc >>
rect 49 539 95 585
rect 263 569 309 615
rect 665 549 711 595
rect 1075 588 1121 634
rect 1322 515 1368 561
rect 1529 670 1575 716
rect 2649 689 2695 735
rect 1777 513 1823 559
rect 1921 525 1967 571
rect 2160 516 2206 562
rect 2897 529 2943 575
rect 3105 582 3151 628
rect 3302 520 3348 566
rect 3506 537 3552 583
rect 3710 516 3756 562
rect 3905 593 3951 639
rect 4111 540 4157 586
rect 4329 593 4375 639
rect 4555 544 4601 590
rect 4703 525 4749 665
rect 4907 525 4953 665
<< polysilicon >>
rect 124 720 988 760
rect 124 628 224 720
rect 348 628 448 672
rect 496 628 596 672
rect 740 628 840 672
rect 888 628 988 720
rect 1185 687 1285 731
rect 1648 720 2336 760
rect 1648 660 1748 720
rect 2236 678 2336 720
rect 124 432 224 502
rect 124 351 244 432
rect 124 305 150 351
rect 196 305 244 351
rect 124 228 244 305
rect 348 351 448 502
rect 496 469 596 502
rect 496 423 525 469
rect 571 423 596 469
rect 496 410 596 423
rect 348 305 374 351
rect 420 305 448 351
rect 348 272 448 305
rect 740 407 840 502
rect 888 458 988 502
rect 740 361 753 407
rect 799 361 840 407
rect 1185 415 1285 502
rect 1996 622 2096 666
rect 2236 632 2264 678
rect 2310 632 2336 678
rect 2476 641 2576 685
rect 2976 720 4082 760
rect 2768 641 2868 685
rect 2976 641 3076 720
rect 2236 599 2336 632
rect 1185 369 1213 415
rect 1259 413 1285 415
rect 1648 448 1748 497
rect 1259 369 1305 413
rect 740 272 840 361
rect 908 335 1028 363
rect 908 289 926 335
rect 972 289 1028 335
rect 348 228 468 272
rect 516 228 636 272
rect 740 228 860 272
rect 908 228 1028 289
rect 1185 228 1305 369
rect 1648 402 1661 448
rect 1707 402 1748 448
rect 1648 277 1748 402
rect 1996 407 2096 497
rect 3377 628 3477 672
rect 3581 628 3681 672
rect 3982 652 4082 720
rect 4426 712 4526 756
rect 4778 716 4878 760
rect 4186 652 4286 696
rect 2236 430 2336 474
rect 2476 430 2576 516
rect 1996 361 2009 407
rect 2055 376 2096 407
rect 2488 384 2576 430
rect 2768 459 2868 516
rect 2768 413 2794 459
rect 2840 413 2868 459
rect 2768 400 2868 413
rect 2055 361 2404 376
rect 1996 336 2404 361
rect 2284 324 2404 336
rect 2284 278 2325 324
rect 2371 278 2404 324
rect 124 64 244 156
rect 348 112 468 156
rect 516 64 636 156
rect 740 112 860 156
rect 908 112 1028 156
rect 1648 232 1768 277
rect 2060 196 2180 240
rect 2284 196 2404 278
rect 2488 367 2608 384
rect 2488 321 2526 367
rect 2572 321 2608 367
rect 2488 196 2608 321
rect 2788 301 2868 400
rect 2976 301 3076 516
rect 3377 470 3477 503
rect 3377 424 3404 470
rect 3450 424 3477 470
rect 3377 357 3477 424
rect 3581 389 3681 503
rect 3982 451 4082 527
rect 3885 393 4082 451
rect 4186 419 4286 527
rect 3581 363 3766 389
rect 2788 257 2908 301
rect 2956 257 3076 301
rect 3180 336 3300 349
rect 3180 290 3218 336
rect 3264 290 3300 336
rect 3377 317 3524 357
rect 3581 317 3707 363
rect 3753 317 3766 363
rect 3180 257 3300 290
rect 3404 257 3524 317
rect 3650 304 3766 317
rect 3885 377 4005 393
rect 3885 331 3931 377
rect 3977 331 4005 377
rect 4186 373 4223 419
rect 4269 373 4286 419
rect 4186 345 4286 373
rect 1185 91 1305 135
rect 124 24 636 64
rect 1648 64 1768 139
rect 2788 141 2908 185
rect 2956 141 3076 185
rect 3180 141 3300 185
rect 3404 141 3524 185
rect 3885 178 4005 331
rect 4110 305 4286 345
rect 4426 438 4526 527
rect 4426 392 4449 438
rect 4495 392 4526 438
rect 4426 332 4526 392
rect 4778 358 4878 472
rect 4110 178 4230 305
rect 4370 292 4526 332
rect 4738 345 4878 358
rect 4738 299 4752 345
rect 4798 299 4878 345
rect 4738 292 4878 299
rect 4370 199 4490 292
rect 4738 232 4858 292
rect 2060 64 2180 124
rect 2284 80 2404 124
rect 2488 80 2608 124
rect 1648 24 2180 64
rect 3885 62 4005 106
rect 4110 62 4230 106
rect 4370 62 4490 106
rect 4738 24 4858 68
<< polycontact >>
rect 150 305 196 351
rect 525 423 571 469
rect 374 305 420 351
rect 753 361 799 407
rect 2264 632 2310 678
rect 1213 369 1259 415
rect 926 289 972 335
rect 1661 402 1707 448
rect 2009 361 2055 407
rect 2794 413 2840 459
rect 2325 278 2371 324
rect 2526 321 2572 367
rect 3404 424 3450 470
rect 3218 290 3264 336
rect 3707 317 3753 363
rect 3931 331 3977 377
rect 4223 373 4269 419
rect 4449 392 4495 438
rect 4752 299 4798 345
<< metal1 >>
rect 0 735 5040 844
rect 0 724 2649 735
rect 252 615 320 724
rect 49 585 95 608
rect 252 569 263 615
rect 309 569 320 615
rect 1075 634 1121 724
rect 1518 716 1586 724
rect 654 549 665 595
rect 711 549 824 595
rect 1075 577 1121 588
rect 1217 632 1472 678
rect 1518 670 1529 716
rect 1575 670 1586 716
rect 2638 689 2649 724
rect 2695 724 5040 735
rect 2695 689 2706 724
rect 49 523 95 539
rect 778 531 824 549
rect 1217 531 1263 632
rect 1426 624 1472 632
rect 1641 632 1967 678
rect 2253 632 2264 678
rect 2310 643 2556 678
rect 2752 643 3046 678
rect 2310 632 3046 643
rect 1641 624 1687 632
rect 1426 578 1687 624
rect 49 477 571 523
rect 778 484 1263 531
rect 1322 561 1368 578
rect 1777 559 1823 578
rect 1368 515 1707 524
rect 1322 477 1707 515
rect 49 215 95 477
rect 525 469 571 477
rect 49 156 95 169
rect 141 351 206 430
rect 141 305 150 351
rect 196 305 206 351
rect 141 119 206 305
rect 365 351 430 430
rect 365 305 374 351
rect 420 305 430 351
rect 273 215 319 228
rect 273 60 319 169
rect 365 119 430 305
rect 525 307 571 423
rect 682 407 878 431
rect 682 361 753 407
rect 799 361 878 407
rect 682 353 878 361
rect 1026 415 1326 431
rect 1026 369 1213 415
rect 1259 369 1326 415
rect 1026 353 1326 369
rect 926 335 972 348
rect 525 289 926 307
rect 525 261 972 289
rect 1018 252 1248 298
rect 1389 255 1435 477
rect 1661 448 1707 477
rect 1661 382 1707 402
rect 1777 407 1823 513
rect 1921 571 1967 632
rect 2510 597 2798 632
rect 2897 575 2943 586
rect 1921 497 1967 525
rect 2160 562 2206 574
rect 2160 459 2206 516
rect 2160 413 2794 459
rect 2840 413 2851 459
rect 2897 444 2943 529
rect 3000 536 3046 632
rect 3092 628 3164 724
rect 3092 582 3105 628
rect 3151 582 3164 628
rect 3210 623 3450 669
rect 3210 536 3256 623
rect 3000 490 3256 536
rect 3302 566 3348 577
rect 3302 444 3348 520
rect 1777 361 2009 407
rect 2055 361 2078 407
rect 1777 360 2078 361
rect 1018 215 1064 252
rect 650 169 665 215
rect 711 169 1064 215
rect 1110 194 1156 205
rect 1110 60 1156 148
rect 1202 152 1248 252
rect 1367 244 1435 255
rect 1367 198 1378 244
rect 1424 198 1435 244
rect 1481 259 1736 306
rect 1481 152 1527 259
rect 1202 106 1527 152
rect 1573 198 1619 209
rect 1573 60 1619 152
rect 1690 152 1736 259
rect 1830 244 1898 360
rect 1830 198 1841 244
rect 1887 198 1898 244
rect 1985 183 2031 196
rect 1690 137 1985 152
rect 1690 106 2031 137
rect 2209 183 2255 413
rect 2897 398 3348 444
rect 3404 470 3450 623
rect 3404 413 3450 424
rect 3506 623 3848 669
rect 3506 583 3552 623
rect 2897 367 2943 398
rect 2325 324 2391 340
rect 2371 278 2391 324
rect 2495 321 2526 367
rect 2572 321 2943 367
rect 2325 275 2391 278
rect 2325 229 2866 275
rect 2209 124 2255 137
rect 2624 137 2637 183
rect 2683 137 2696 183
rect 2624 60 2696 137
rect 2820 152 2866 229
rect 3094 244 3162 398
rect 3506 352 3552 537
rect 3710 562 3756 577
rect 3710 463 3756 516
rect 3802 547 3848 623
rect 3894 639 3962 724
rect 3894 593 3905 639
rect 3951 593 3962 639
rect 4008 632 4268 678
rect 4008 547 4054 632
rect 3802 501 4054 547
rect 4100 540 4111 586
rect 4157 540 4168 586
rect 3094 198 3105 244
rect 3151 198 3162 244
rect 3218 336 3264 348
rect 3218 152 3264 290
rect 3318 305 3552 352
rect 3598 455 3756 463
rect 3598 409 3856 455
rect 3318 244 3386 305
rect 3598 253 3644 409
rect 3318 198 3329 244
rect 3375 198 3386 244
rect 3542 244 3644 253
rect 3542 198 3553 244
rect 3599 198 3644 244
rect 3690 317 3707 363
rect 3753 317 3764 363
rect 3690 152 3764 317
rect 2820 106 3764 152
rect 3810 165 3856 409
rect 3924 377 4022 438
rect 3924 331 3931 377
rect 3977 331 4022 377
rect 3924 234 4022 331
rect 4100 152 4168 540
rect 4222 547 4268 632
rect 4318 639 4386 724
rect 4318 593 4329 639
rect 4375 593 4386 639
rect 4703 665 4749 724
rect 4555 590 4601 630
rect 4222 501 4506 547
rect 4438 438 4506 501
rect 4223 419 4269 434
rect 4438 392 4449 438
rect 4495 392 4506 438
rect 4223 345 4269 373
rect 4555 356 4601 544
rect 4703 506 4749 525
rect 4844 665 4954 676
rect 4844 525 4907 665
rect 4953 525 4954 665
rect 4555 345 4798 356
rect 4223 299 4752 345
rect 4508 288 4798 299
rect 4508 186 4578 288
rect 3856 119 4168 152
rect 3810 106 4168 119
rect 4295 165 4341 178
rect 4508 140 4519 186
rect 4565 140 4578 186
rect 4508 131 4578 140
rect 4663 142 4709 181
rect 4295 60 4341 119
rect 4844 177 4954 525
rect 4844 131 4887 177
rect 4933 131 4954 177
rect 4844 119 4954 131
rect 4663 60 4709 96
rect 0 -60 5040 60
<< labels >>
flabel metal1 s 4844 119 4954 676 0 FreeSans 400 0 0 0 Q
port 6 nsew default output
flabel metal1 s 141 119 206 430 0 FreeSans 400 0 0 0 SE
port 2 nsew default input
flabel metal1 s 3924 234 4022 438 0 FreeSans 400 0 0 0 SETN
port 3 nsew default input
flabel metal1 s 365 119 430 430 0 FreeSans 400 0 0 0 SI
port 4 nsew default input
flabel metal1 s 0 724 5040 844 0 FreeSans 400 0 0 0 VDD
port 7 nsew power bidirectional abutment
flabel metal1 s 273 209 319 228 0 FreeSans 400 0 0 0 VSS
port 10 nsew ground bidirectional abutment
flabel metal1 s 1026 353 1326 431 0 FreeSans 400 0 0 0 CLK
port 5 nsew clock input
flabel metal1 s 682 353 878 431 0 FreeSans 400 0 0 0 D
port 1 nsew default input
flabel nwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_mcu_sc7
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v1
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 4703 689 4749 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4318 689 4386 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3894 689 3962 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3092 689 3164 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2638 689 2706 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1518 689 1586 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 689 1121 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 689 320 724 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 670 4749 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4318 670 4386 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3894 670 3962 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3092 670 3164 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1518 670 1586 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 670 1121 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 670 320 689 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 593 4749 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4318 593 4386 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3894 593 3962 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3092 593 3164 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 593 1121 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 593 320 670 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 582 4749 593 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 3092 582 3164 593 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 582 1121 593 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 582 320 593 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 577 4749 582 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1075 577 1121 582 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 577 320 582 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 569 4749 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 252 569 320 577 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 4703 506 4749 569 1 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1573 205 1619 209 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 205 319 209 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1573 183 1619 205 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1110 183 1156 205 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 183 319 205 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2624 181 2696 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1573 181 1619 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1110 181 1156 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 181 319 183 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4663 178 4709 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2624 178 2696 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1573 178 1619 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1110 178 1156 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 178 319 181 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4663 60 4709 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 4295 60 4341 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 2624 60 2696 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1573 60 1619 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 1110 60 1156 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 60 319 178 1 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 5040 60 1 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 5040 784
string GDS_END 286858
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 275946
string LEFclass core
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
<< end >>
