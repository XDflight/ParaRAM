magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 918 2464 1098
rect 69 775 115 918
rect 731 729 777 871
rect 1373 775 1419 918
rect 1831 729 1877 868
rect 2269 775 2315 918
rect 731 683 2291 729
rect 142 588 1182 634
rect 142 443 203 588
rect 388 454 538 500
rect 584 454 652 542
rect 1136 500 1182 588
rect 1486 588 2199 634
rect 926 454 1090 500
rect 1136 454 1314 500
rect 492 408 538 454
rect 926 408 978 454
rect 1486 443 1547 588
rect 1703 443 1762 542
rect 2153 443 2199 588
rect 492 362 978 408
rect 2245 397 2291 683
rect 926 354 978 362
rect 1598 351 2291 397
rect 273 90 319 219
rect 721 90 767 219
rect 1169 90 1215 219
rect 1598 228 1663 351
rect 2065 228 2111 351
rect 0 -90 2464 90
<< obsm1 >>
rect 49 308 895 313
rect 1011 308 1439 313
rect 49 267 1439 308
rect 49 151 95 267
rect 497 151 543 267
rect 874 262 1032 267
rect 945 146 1032 262
rect 1393 182 1439 267
rect 1841 182 1887 305
rect 2337 182 2383 313
rect 1393 136 2383 182
<< labels >>
rlabel metal1 s 584 454 652 542 6 A1
port 1 nsew default input
rlabel metal1 s 926 454 1090 500 6 A2
port 2 nsew default input
rlabel metal1 s 388 454 538 500 6 A2
port 2 nsew default input
rlabel metal1 s 926 408 978 454 6 A2
port 2 nsew default input
rlabel metal1 s 492 408 538 454 6 A2
port 2 nsew default input
rlabel metal1 s 492 362 978 408 6 A2
port 2 nsew default input
rlabel metal1 s 926 354 978 362 6 A2
port 2 nsew default input
rlabel metal1 s 142 588 1182 634 6 A3
port 3 nsew default input
rlabel metal1 s 1136 500 1182 588 6 A3
port 3 nsew default input
rlabel metal1 s 142 500 203 588 6 A3
port 3 nsew default input
rlabel metal1 s 1136 454 1314 500 6 A3
port 3 nsew default input
rlabel metal1 s 142 454 203 500 6 A3
port 3 nsew default input
rlabel metal1 s 142 443 203 454 6 A3
port 3 nsew default input
rlabel metal1 s 1703 443 1762 542 6 B1
port 4 nsew default input
rlabel metal1 s 1486 588 2199 634 6 B2
port 5 nsew default input
rlabel metal1 s 2153 443 2199 588 6 B2
port 5 nsew default input
rlabel metal1 s 1486 443 1547 588 6 B2
port 5 nsew default input
rlabel metal1 s 731 868 777 871 6 ZN
port 6 nsew default output
rlabel metal1 s 1831 729 1877 868 6 ZN
port 6 nsew default output
rlabel metal1 s 731 729 777 868 6 ZN
port 6 nsew default output
rlabel metal1 s 731 683 2291 729 6 ZN
port 6 nsew default output
rlabel metal1 s 2245 397 2291 683 6 ZN
port 6 nsew default output
rlabel metal1 s 1598 351 2291 397 6 ZN
port 6 nsew default output
rlabel metal1 s 2065 228 2111 351 6 ZN
port 6 nsew default output
rlabel metal1 s 1598 228 1663 351 6 ZN
port 6 nsew default output
rlabel metal1 s 0 918 2464 1098 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 2269 775 2315 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1373 775 1419 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 69 775 115 918 6 VDD
port 7 nsew power bidirectional abutment
rlabel metal1 s 1169 90 1215 219 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 721 90 767 219 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 273 90 319 219 6 VSS
port 8 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 2464 90 8 VSS
port 8 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2464 1008
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 167966
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 162240
<< end >>
