magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 120 1474
rect 224 0 344 1474
rect 448 0 568 1474
rect 672 0 792 1474
rect 896 0 1016 1474
rect 1120 0 1240 1474
rect 1344 0 1464 1474
rect 1568 0 1688 1474
rect 1792 0 1912 1474
rect 2016 0 2136 1474
rect 2240 0 2360 1474
rect 2464 0 2584 1474
rect 2688 0 2808 1474
rect 2912 0 3032 1474
rect 3136 0 3256 1474
rect 3360 0 3480 1474
rect 3584 0 3704 1474
rect 3808 0 3928 1474
rect 4032 0 4152 1474
rect 4256 0 4376 1474
<< mvndiff >>
rect -88 1461 0 1474
rect -88 13 -75 1461
rect -29 13 0 1461
rect -88 0 0 13
rect 120 1461 224 1474
rect 120 13 149 1461
rect 195 13 224 1461
rect 120 0 224 13
rect 344 1461 448 1474
rect 344 13 373 1461
rect 419 13 448 1461
rect 344 0 448 13
rect 568 1461 672 1474
rect 568 13 597 1461
rect 643 13 672 1461
rect 568 0 672 13
rect 792 1461 896 1474
rect 792 13 821 1461
rect 867 13 896 1461
rect 792 0 896 13
rect 1016 1461 1120 1474
rect 1016 13 1045 1461
rect 1091 13 1120 1461
rect 1016 0 1120 13
rect 1240 1461 1344 1474
rect 1240 13 1269 1461
rect 1315 13 1344 1461
rect 1240 0 1344 13
rect 1464 1461 1568 1474
rect 1464 13 1493 1461
rect 1539 13 1568 1461
rect 1464 0 1568 13
rect 1688 1461 1792 1474
rect 1688 13 1717 1461
rect 1763 13 1792 1461
rect 1688 0 1792 13
rect 1912 1461 2016 1474
rect 1912 13 1941 1461
rect 1987 13 2016 1461
rect 1912 0 2016 13
rect 2136 1461 2240 1474
rect 2136 13 2165 1461
rect 2211 13 2240 1461
rect 2136 0 2240 13
rect 2360 1461 2464 1474
rect 2360 13 2389 1461
rect 2435 13 2464 1461
rect 2360 0 2464 13
rect 2584 1461 2688 1474
rect 2584 13 2613 1461
rect 2659 13 2688 1461
rect 2584 0 2688 13
rect 2808 1461 2912 1474
rect 2808 13 2837 1461
rect 2883 13 2912 1461
rect 2808 0 2912 13
rect 3032 1461 3136 1474
rect 3032 13 3061 1461
rect 3107 13 3136 1461
rect 3032 0 3136 13
rect 3256 1461 3360 1474
rect 3256 13 3285 1461
rect 3331 13 3360 1461
rect 3256 0 3360 13
rect 3480 1461 3584 1474
rect 3480 13 3509 1461
rect 3555 13 3584 1461
rect 3480 0 3584 13
rect 3704 1461 3808 1474
rect 3704 13 3733 1461
rect 3779 13 3808 1461
rect 3704 0 3808 13
rect 3928 1461 4032 1474
rect 3928 13 3957 1461
rect 4003 13 4032 1461
rect 3928 0 4032 13
rect 4152 1461 4256 1474
rect 4152 13 4181 1461
rect 4227 13 4256 1461
rect 4152 0 4256 13
rect 4376 1461 4464 1474
rect 4376 13 4405 1461
rect 4451 13 4464 1461
rect 4376 0 4464 13
<< mvndiffc >>
rect -75 13 -29 1461
rect 149 13 195 1461
rect 373 13 419 1461
rect 597 13 643 1461
rect 821 13 867 1461
rect 1045 13 1091 1461
rect 1269 13 1315 1461
rect 1493 13 1539 1461
rect 1717 13 1763 1461
rect 1941 13 1987 1461
rect 2165 13 2211 1461
rect 2389 13 2435 1461
rect 2613 13 2659 1461
rect 2837 13 2883 1461
rect 3061 13 3107 1461
rect 3285 13 3331 1461
rect 3509 13 3555 1461
rect 3733 13 3779 1461
rect 3957 13 4003 1461
rect 4181 13 4227 1461
rect 4405 13 4451 1461
<< polysilicon >>
rect 0 1474 120 1518
rect 224 1474 344 1518
rect 448 1474 568 1518
rect 672 1474 792 1518
rect 896 1474 1016 1518
rect 1120 1474 1240 1518
rect 1344 1474 1464 1518
rect 1568 1474 1688 1518
rect 1792 1474 1912 1518
rect 2016 1474 2136 1518
rect 2240 1474 2360 1518
rect 2464 1474 2584 1518
rect 2688 1474 2808 1518
rect 2912 1474 3032 1518
rect 3136 1474 3256 1518
rect 3360 1474 3480 1518
rect 3584 1474 3704 1518
rect 3808 1474 3928 1518
rect 4032 1474 4152 1518
rect 4256 1474 4376 1518
rect 0 -44 120 0
rect 224 -44 344 0
rect 448 -44 568 0
rect 672 -44 792 0
rect 896 -44 1016 0
rect 1120 -44 1240 0
rect 1344 -44 1464 0
rect 1568 -44 1688 0
rect 1792 -44 1912 0
rect 2016 -44 2136 0
rect 2240 -44 2360 0
rect 2464 -44 2584 0
rect 2688 -44 2808 0
rect 2912 -44 3032 0
rect 3136 -44 3256 0
rect 3360 -44 3480 0
rect 3584 -44 3704 0
rect 3808 -44 3928 0
rect 4032 -44 4152 0
rect 4256 -44 4376 0
<< metal1 >>
rect -75 1461 -29 1474
rect -75 0 -29 13
rect 149 1461 195 1474
rect 149 0 195 13
rect 373 1461 419 1474
rect 373 0 419 13
rect 597 1461 643 1474
rect 597 0 643 13
rect 821 1461 867 1474
rect 821 0 867 13
rect 1045 1461 1091 1474
rect 1045 0 1091 13
rect 1269 1461 1315 1474
rect 1269 0 1315 13
rect 1493 1461 1539 1474
rect 1493 0 1539 13
rect 1717 1461 1763 1474
rect 1717 0 1763 13
rect 1941 1461 1987 1474
rect 1941 0 1987 13
rect 2165 1461 2211 1474
rect 2165 0 2211 13
rect 2389 1461 2435 1474
rect 2389 0 2435 13
rect 2613 1461 2659 1474
rect 2613 0 2659 13
rect 2837 1461 2883 1474
rect 2837 0 2883 13
rect 3061 1461 3107 1474
rect 3061 0 3107 13
rect 3285 1461 3331 1474
rect 3285 0 3331 13
rect 3509 1461 3555 1474
rect 3509 0 3555 13
rect 3733 1461 3779 1474
rect 3733 0 3779 13
rect 3957 1461 4003 1474
rect 3957 0 4003 13
rect 4181 1461 4227 1474
rect 4181 0 4227 13
rect 4405 1461 4451 1474
rect 4405 0 4451 13
<< labels >>
flabel metal1 s -52 737 -52 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 4428 737 4428 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 172 737 172 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 396 737 396 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 620 737 620 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 844 737 844 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 1068 737 1068 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 1292 737 1292 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 1516 737 1516 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 1740 737 1740 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 1964 737 1964 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 2188 737 2188 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 2412 737 2412 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 2636 737 2636 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 2860 737 2860 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 3084 737 3084 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 3308 737 3308 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 3532 737 3532 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 3756 737 3756 737 0 FreeSans 200 0 0 0 D
flabel metal1 s 3980 737 3980 737 0 FreeSans 200 0 0 0 S
flabel metal1 s 4204 737 4204 737 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 498206
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 471172
<< end >>
