magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -203 10266 787 12370
rect -7 8752 622 10266
rect -7 8695 624 8752
rect -5 7108 624 8695
rect -221 1164 756 1620
rect -203 648 756 1164
<< pmos >>
rect 102 11191 222 11873
rect 327 11191 447 11873
rect 102 10416 222 11098
rect 327 10416 447 11098
rect 67 788 187 1085
rect 318 788 438 1085
<< pdiff >>
rect -4 11191 102 11873
rect 222 11191 327 11873
rect 447 11191 553 11873
rect -4 10416 102 11098
rect 222 10416 327 11098
rect 447 10416 553 11098
rect -67 960 67 1085
rect -67 914 -23 960
rect 23 914 67 960
rect -67 788 67 914
rect 187 960 318 1085
rect 187 914 230 960
rect 276 914 318 960
rect 187 788 318 914
rect 438 960 620 1085
rect 438 914 480 960
rect 526 914 620 960
rect 438 788 620 914
<< pdiffc >>
rect -23 914 23 960
rect 230 914 276 960
rect 480 914 526 960
<< psubdiff >>
rect -80 5260 80 5320
rect -80 5214 -23 5260
rect 23 5214 80 5260
rect -80 5154 80 5214
rect 540 5260 700 5320
rect 540 5214 597 5260
rect 643 5214 700 5260
rect 540 5154 700 5214
rect -80 96 620 155
rect -80 50 -23 96
rect 23 50 135 96
rect 181 50 293 96
rect 339 50 451 96
rect 497 50 620 96
rect -80 -10 620 50
<< nsubdiff >>
rect -1 12165 651 12222
rect -1 12119 129 12165
rect 175 12119 287 12165
rect 333 12119 445 12165
rect 491 12119 651 12165
rect -1 12062 651 12119
rect -78 1415 620 1472
rect -78 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -78 1312 620 1369
<< psubdiffcont >>
rect -23 5214 23 5260
rect 597 5214 643 5260
rect -23 50 23 96
rect 135 50 181 96
rect 293 50 339 96
rect 451 50 497 96
<< nsubdiffcont >>
rect 129 12119 175 12165
rect 287 12119 333 12165
rect 445 12119 491 12165
rect -23 1369 23 1415
rect 135 1369 181 1415
rect 293 1369 339 1415
rect 451 1369 497 1415
<< polysilicon >>
rect 102 11873 222 11946
rect 327 11873 447 11946
rect 102 11098 222 11191
rect 327 11098 447 11191
rect 102 10348 222 10416
rect 327 10348 447 10416
rect 102 10329 447 10348
rect 102 10283 155 10329
rect 389 10283 447 10329
rect 102 10264 447 10283
rect 248 10198 368 10264
rect 248 8764 368 8836
rect 250 8611 370 8684
rect 250 7164 370 7249
rect 250 7118 293 7164
rect 339 7118 370 7164
rect 250 7099 370 7118
rect 250 4930 370 5505
rect 250 3469 370 3520
rect 250 3423 287 3469
rect 333 3423 370 3469
rect 250 3404 370 3423
rect 250 3192 370 3211
rect 250 3146 287 3192
rect 333 3146 370 3192
rect 250 3095 370 3146
rect 67 1225 438 1244
rect 67 1179 230 1225
rect 276 1179 438 1225
rect 67 1145 438 1179
rect 67 1085 187 1145
rect 318 1085 438 1145
rect 67 635 187 788
rect 318 636 438 788
rect 52 598 187 635
rect 276 602 438 636
rect 52 539 172 598
rect 276 539 396 602
rect 52 497 170 498
rect 52 310 172 382
rect 276 310 396 382
<< polycontact >>
rect 155 10283 389 10329
rect 293 7118 339 7164
rect 287 3423 333 3469
rect 287 3146 333 3192
rect 230 1179 276 1225
<< metal1 >>
rect -58 12203 620 12227
rect -58 12165 281 12203
rect 333 12165 620 12203
rect -58 12119 129 12165
rect 175 12151 281 12165
rect 175 12119 287 12151
rect 333 12119 445 12165
rect 491 12119 620 12165
rect -58 12017 620 12119
rect -58 11965 281 12017
rect 333 11965 620 12017
rect -58 11944 620 11965
rect -58 10425 58 11944
rect 217 11633 333 11864
rect 217 11581 259 11633
rect 311 11581 333 11633
rect 217 11447 333 11581
rect 217 11395 259 11447
rect 311 11395 333 11447
rect 217 11200 333 11395
rect 217 10858 333 11089
rect 217 10702 249 10858
rect 301 10702 333 10858
rect 217 10425 333 10702
rect 478 10425 620 11944
rect 144 10329 400 10340
rect 144 10283 155 10329
rect 389 10283 400 10329
rect 144 10272 400 10283
rect 62 9638 219 9650
rect 62 9482 74 9638
rect 126 9482 219 9638
rect 62 9470 219 9482
rect 397 9638 556 9650
rect 397 9482 492 9638
rect 544 9482 556 9638
rect 397 9470 556 9482
rect 74 8598 192 8610
rect 74 8442 86 8598
rect 138 8442 192 8598
rect 74 8045 192 8442
rect 114 7525 192 8045
rect 74 7248 192 7525
rect 434 7248 550 8602
rect 74 6919 162 7248
rect 219 7166 401 7178
rect 219 7010 290 7166
rect 342 7010 401 7166
rect 219 6995 401 7010
rect 458 6919 550 7248
rect 74 5567 192 6919
rect 434 5657 550 6919
rect 399 5567 550 5657
rect 399 5487 445 5567
rect 45 5465 445 5487
rect 45 5413 75 5465
rect 127 5413 445 5465
rect 45 5390 445 5413
rect -71 5306 71 5311
rect 549 5306 691 5311
rect -71 5267 691 5306
rect -71 5260 347 5267
rect -71 5214 -23 5260
rect 23 5215 347 5260
rect 399 5260 691 5267
rect 399 5215 597 5260
rect 23 5214 597 5215
rect 643 5214 691 5260
rect -71 5172 691 5214
rect -71 5163 71 5172
rect 549 5163 691 5172
rect 48 5058 561 5084
rect 48 5006 492 5058
rect 544 5006 561 5058
rect 48 4987 561 5006
rect 48 3553 188 4987
rect 431 3553 550 4907
rect 48 3060 145 3553
rect 219 3469 401 3483
rect 219 3459 287 3469
rect 333 3459 401 3469
rect 219 3407 286 3459
rect 338 3407 401 3459
rect 219 3348 401 3407
rect 219 3196 401 3268
rect 219 3144 284 3196
rect 336 3144 401 3196
rect 219 3132 401 3144
rect 464 3060 550 3553
rect 48 1708 188 3060
rect 431 1710 550 3060
rect 421 1554 550 1710
rect -58 1415 620 1452
rect -58 1369 -23 1415
rect 23 1369 135 1415
rect 181 1369 293 1415
rect 339 1369 451 1415
rect 497 1369 620 1415
rect -58 1332 620 1369
rect -58 960 58 1332
rect 136 1228 405 1252
rect 136 1225 287 1228
rect 136 1179 230 1225
rect 276 1179 287 1225
rect 136 1176 287 1179
rect 339 1176 405 1228
rect 136 1155 405 1176
rect 548 1076 620 1332
rect -58 914 -23 960
rect 23 914 58 960
rect -58 797 58 914
rect 195 1064 324 1076
rect 195 908 207 1064
rect 259 960 324 1064
rect 276 914 324 960
rect 259 908 324 914
rect 195 797 324 908
rect 445 960 620 1076
rect 445 914 480 960
rect 526 914 620 960
rect 445 797 620 914
rect 217 500 289 797
rect -58 271 58 500
rect 192 380 289 500
rect 425 271 620 500
rect -58 147 620 271
rect -71 96 620 147
rect -71 50 -23 96
rect 23 50 135 96
rect 181 50 293 96
rect 339 50 451 96
rect 497 50 620 96
rect -71 -1 620 50
<< via1 >>
rect 281 12165 333 12203
rect 281 12151 287 12165
rect 287 12151 333 12165
rect 281 11965 333 12017
rect 259 11581 311 11633
rect 259 11395 311 11447
rect 249 10702 301 10858
rect 74 9482 126 9638
rect 492 9482 544 9638
rect 86 8442 138 8598
rect 290 7164 342 7166
rect 290 7118 293 7164
rect 293 7118 339 7164
rect 339 7118 342 7164
rect 290 7010 342 7118
rect 75 5413 127 5465
rect 347 5215 399 5267
rect 492 5006 544 5058
rect 286 3423 287 3459
rect 287 3423 333 3459
rect 333 3423 338 3459
rect 286 3407 338 3423
rect 284 3192 336 3196
rect 284 3146 287 3192
rect 287 3146 333 3192
rect 333 3146 336 3192
rect 284 3144 336 3146
rect 287 1176 339 1228
rect 207 960 259 1064
rect 207 914 230 960
rect 230 914 259 960
rect 207 908 259 914
<< metal2 >>
rect 72 11584 128 12275
rect 245 12205 374 12227
rect 245 12149 279 12205
rect 335 12149 374 12205
rect 245 12019 374 12149
rect 245 11963 279 12019
rect 335 11963 374 12019
rect 245 11944 374 11963
rect 239 11633 331 11673
rect 239 11584 259 11633
rect 72 11581 259 11584
rect 311 11581 331 11633
rect 72 11528 331 11581
rect 72 9650 128 11528
rect 239 11447 331 11528
rect 239 11395 259 11447
rect 311 11395 331 11447
rect 239 11355 331 11395
rect 237 10858 313 10870
rect 237 10702 249 10858
rect 301 10808 313 10858
rect 490 10808 546 12275
rect 301 10752 546 10808
rect 301 10702 313 10752
rect 237 10690 313 10702
rect 490 9650 546 10752
rect 62 9638 138 9650
rect 62 9482 74 9638
rect 126 9482 138 9638
rect 62 9470 138 9482
rect 480 9638 556 9650
rect 480 9482 492 9638
rect 544 9482 556 9638
rect 480 9470 556 9482
rect 72 8610 128 9470
rect 72 8598 150 8610
rect 72 8442 86 8598
rect 138 8442 150 8598
rect 72 8430 150 8442
rect 278 7166 354 7178
rect 278 7010 290 7166
rect 342 7010 354 7166
rect 278 6998 354 7010
rect 0 5465 139 5477
rect 0 5413 75 5465
rect 127 5413 139 5465
rect 0 5401 139 5413
rect 288 5397 344 6998
rect 199 5341 344 5397
rect 199 3655 255 5341
rect 335 5267 411 5279
rect 335 5256 347 5267
rect 399 5256 411 5267
rect 335 5096 345 5256
rect 401 5096 411 5256
rect 335 5086 411 5096
rect 490 5070 546 9470
rect 480 5058 556 5070
rect 480 5006 492 5058
rect 544 5006 556 5058
rect 480 4994 556 5006
rect 113 3599 255 3655
rect 113 3197 169 3599
rect 480 3483 574 4517
rect 250 3459 574 3483
rect 250 3407 286 3459
rect 338 3407 574 3459
rect 250 3386 574 3407
rect 272 3197 348 3208
rect 113 3196 348 3197
rect 113 3144 284 3196
rect 336 3144 348 3196
rect 113 3141 348 3144
rect 113 1076 169 3141
rect 272 3132 348 3141
rect 480 1853 574 3386
rect 275 1756 574 1853
rect 275 1228 351 1756
rect 275 1176 287 1228
rect 339 1176 351 1228
rect 275 1155 351 1176
rect 113 1064 271 1076
rect 113 908 207 1064
rect 259 908 271 1064
rect 113 896 271 908
rect 245 49 374 278
<< via2 >>
rect 279 12203 335 12205
rect 279 12151 281 12203
rect 281 12151 333 12203
rect 333 12151 335 12203
rect 279 12149 335 12151
rect 279 12017 335 12019
rect 279 11965 281 12017
rect 281 11965 333 12017
rect 333 11965 335 12017
rect 279 11963 335 11965
rect 345 5215 347 5256
rect 347 5215 399 5256
rect 399 5215 401 5256
rect 345 5096 401 5215
<< metal3 >>
rect -65 12205 651 12347
rect -65 12149 279 12205
rect 335 12149 651 12205
rect -65 12019 651 12149
rect -65 11963 279 12019
rect 335 11963 651 12019
rect -65 10538 651 11963
rect -1 5256 636 6638
rect -1 5096 345 5256
rect 401 5096 636 5256
rect -1 4656 636 5096
rect -1 4331 636 4546
rect -1 4009 636 4224
rect -1 3688 636 3903
rect -1 3366 636 3581
rect -1 2674 636 2889
rect -1 2352 636 2567
rect -1 2030 636 2245
rect -1 1708 636 1923
rect -1 1160 636 1602
rect -1 49 636 504
use M1_NWELL$$46277676_128x8m81  M1_NWELL$$46277676_128x8m81_0
timestamp 1666464484
transform 1 0 310 0 1 12142
box 0 0 1 1
use M1_NWELL$$47121452_128x8m81  M1_NWELL$$47121452_128x8m81_0
timestamp 1666464484
transform 1 0 237 0 1 1392
box 0 0 1 1
use M1_POLY24310590548731_128x8m81  M1_POLY24310590548731_128x8m81_0
timestamp 1666464484
transform 1 0 272 0 1 10306
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_0
timestamp 1666464484
transform 1 0 310 0 1 3446
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_1
timestamp 1666464484
transform 1 0 310 0 1 3169
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_2
timestamp 1666464484
transform 1 0 253 0 1 1202
box 0 0 1 1
use M1_POLY24310590548732_128x8m81  M1_POLY24310590548732_128x8m81_3
timestamp 1666464484
transform 1 0 316 0 1 7141
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_0
timestamp 1666464484
transform 1 0 620 0 1 5237
box 0 0 1 1
use M1_PSUB$$45111340_128x8m81  M1_PSUB$$45111340_128x8m81_1
timestamp 1666464484
transform 1 0 0 0 1 5237
box 0 0 1 1
use M1_PSUB$$47122476_128x8m81  M1_PSUB$$47122476_128x8m81_0
timestamp 1666464484
transform 1 0 237 0 1 73
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_0
timestamp 1666464484
transform 1 0 100 0 1 9560
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_1
timestamp 1666464484
transform 1 0 518 0 1 9560
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_2
timestamp 1666464484
transform 1 0 275 0 1 10780
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_3
timestamp 1666464484
transform 1 0 316 0 1 7088
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_4
timestamp 1666464484
transform 1 0 233 0 1 986
box 0 0 1 1
use M2_M1431059054875_128x8m81  M2_M1431059054875_128x8m81_5
timestamp 1666464484
transform 1 0 112 0 1 8520
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_0
timestamp 1666464484
transform 1 0 373 0 1 5241
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_1
timestamp 1666464484
transform 1 0 518 0 1 5032
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_2
timestamp 1666464484
transform 1 0 313 0 1 1202
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_3
timestamp 1666464484
transform 1 0 310 0 1 3170
box 0 0 1 1
use M2_M14310590548724_128x8m81  M2_M14310590548724_128x8m81_4
timestamp 1666464484
transform 1 0 101 0 1 5439
box 0 0 1 1
use M3_M2431059054871_128x8m81  M3_M2431059054871_128x8m81_0
timestamp 1666464484
transform 1 0 373 0 1 5176
box 0 0 1 1
use nmos_1p2$$47119404_128x8m81  nmos_1p2$$47119404_128x8m81_0
timestamp 1666464484
transform 1 0 281 0 -1 4915
box -119 -74 177 1434
use nmos_1p2$$47119404_128x8m81  nmos_1p2$$47119404_128x8m81_1
timestamp 1666464484
transform 1 0 281 0 -1 6919
box -119 -74 177 1434
use nmos_5p0431059054872_128x8m81  nmos_5p0431059054872_128x8m81_0
timestamp 1666464484
transform 1 0 52 0 1 383
box -88 -44 432 158
use pmos_1p2$$46889004_128x8m81  pmos_1p2$$46889004_128x8m81_0
timestamp 1666464484
transform 1 0 281 0 -1 3060
box -286 -142 343 1502
use pmos_5p0431059054871_128x8m81  pmos_5p0431059054871_128x8m81_0
timestamp 1666464484
transform 1 0 248 0 -1 10197
box -208 -120 328 1482
use pmos_5p0431059054871_128x8m81  pmos_5p0431059054871_128x8m81_1
timestamp 1666464484
transform 1 0 250 0 -1 8610
box -208 -120 328 1482
use via1_2_128x8m81  via1_2_128x8m81_0
timestamp 1666464484
transform 1 0 264 0 1 88
box -1 -1 93 128
use via1_R90_128x8m81  via1_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 378 1 0 3387
box 0 0 1 1
use via1_R90_128x8m81  via1_R90_128x8m81_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
use via1_R90_128x8m81  via1_R90_128x8m81_2
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via1_x2_128x8m81  via1_x2_128x8m81_0
timestamp 1666464484
transform 1 0 239 0 1 11355
box 0 0 1 1
use via2_R90_128x8m81  via2_R90_128x8m81_0
timestamp 1666464484
transform 0 -1 373 1 0 11945
box 0 0 1 1
use via2_R90_128x8m81  via2_R90_128x8m81_1
timestamp 1666464484
transform 0 -1 373 1 0 12131
box 0 0 1 1
<< labels >>
rlabel metal3 s 279 91 279 91 4 vss
port 1 nsew
rlabel metal3 s 318 12094 318 12094 4 vdd
port 2 nsew
rlabel metal3 s 303 5255 303 5255 4 vss
port 1 nsew
rlabel metal2 s 518 11931 518 11931 4 b
port 3 nsew
rlabel metal2 s 105 11931 105 11931 4 bb
port 4 nsew
rlabel metal2 s 0 304 0 304 4 db
port 5 nsew
rlabel metal2 s 285 1222 285 1222 4 ypass
port 6 nsew
rlabel metal1 s 492 1805 492 1805 4 d
port 7 nsew
rlabel metal1 s 259 10272 259 10272 4 pcb
port 8 nsew
rlabel metal1 s 318 1356 318 1356 4 vdd
port 2 nsew
<< properties >>
string GDS_END 198916
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram128x8m8wm1.gds
string GDS_START 189724
string path 1.245 53.900 2.590 53.900 
<< end >>
