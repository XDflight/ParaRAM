magic
tech gf180mcuC
magscale 1 10
timestamp 1666464484
<< metal2 >>
rect -1857 246 1856 284
rect -1857 190 -1820 246
rect -1764 190 -1609 246
rect -1553 190 -1399 246
rect -1343 190 -1188 246
rect -1132 190 -977 246
rect -921 190 -766 246
rect -710 190 -555 246
rect -499 190 -345 246
rect -289 190 -134 246
rect -78 190 78 246
rect 134 190 289 246
rect 345 190 499 246
rect 555 190 710 246
rect 766 190 921 246
rect 977 190 1132 246
rect 1188 190 1343 246
rect 1399 190 1553 246
rect 1609 190 1764 246
rect 1820 190 1856 246
rect -1857 28 1856 190
rect -1857 -28 -1820 28
rect -1764 -28 -1609 28
rect -1553 -28 -1399 28
rect -1343 -28 -1188 28
rect -1132 -28 -977 28
rect -921 -28 -766 28
rect -710 -28 -555 28
rect -499 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 499 28
rect 555 -28 710 28
rect 766 -28 921 28
rect 977 -28 1132 28
rect 1188 -28 1343 28
rect 1399 -28 1553 28
rect 1609 -28 1764 28
rect 1820 -28 1856 28
rect -1857 -190 1856 -28
rect -1857 -246 -1820 -190
rect -1764 -246 -1609 -190
rect -1553 -246 -1399 -190
rect -1343 -246 -1188 -190
rect -1132 -246 -977 -190
rect -921 -246 -766 -190
rect -710 -246 -555 -190
rect -499 -246 -345 -190
rect -289 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 289 -190
rect 345 -246 499 -190
rect 555 -246 710 -190
rect 766 -246 921 -190
rect 977 -246 1132 -190
rect 1188 -246 1343 -190
rect 1399 -246 1553 -190
rect 1609 -246 1764 -190
rect 1820 -246 1856 -190
rect -1857 -284 1856 -246
<< via2 >>
rect -1820 190 -1764 246
rect -1609 190 -1553 246
rect -1399 190 -1343 246
rect -1188 190 -1132 246
rect -977 190 -921 246
rect -766 190 -710 246
rect -555 190 -499 246
rect -345 190 -289 246
rect -134 190 -78 246
rect 78 190 134 246
rect 289 190 345 246
rect 499 190 555 246
rect 710 190 766 246
rect 921 190 977 246
rect 1132 190 1188 246
rect 1343 190 1399 246
rect 1553 190 1609 246
rect 1764 190 1820 246
rect -1820 -28 -1764 28
rect -1609 -28 -1553 28
rect -1399 -28 -1343 28
rect -1188 -28 -1132 28
rect -977 -28 -921 28
rect -766 -28 -710 28
rect -555 -28 -499 28
rect -345 -28 -289 28
rect -134 -28 -78 28
rect 78 -28 134 28
rect 289 -28 345 28
rect 499 -28 555 28
rect 710 -28 766 28
rect 921 -28 977 28
rect 1132 -28 1188 28
rect 1343 -28 1399 28
rect 1553 -28 1609 28
rect 1764 -28 1820 28
rect -1820 -246 -1764 -190
rect -1609 -246 -1553 -190
rect -1399 -246 -1343 -190
rect -1188 -246 -1132 -190
rect -977 -246 -921 -190
rect -766 -246 -710 -190
rect -555 -246 -499 -190
rect -345 -246 -289 -190
rect -134 -246 -78 -190
rect 78 -246 134 -190
rect 289 -246 345 -190
rect 499 -246 555 -190
rect 710 -246 766 -190
rect 921 -246 977 -190
rect 1132 -246 1188 -190
rect 1343 -246 1399 -190
rect 1553 -246 1609 -190
rect 1764 -246 1820 -190
<< metal3 >>
rect -1857 246 1857 284
rect -1857 190 -1820 246
rect -1764 190 -1609 246
rect -1553 190 -1399 246
rect -1343 190 -1188 246
rect -1132 190 -977 246
rect -921 190 -766 246
rect -710 190 -555 246
rect -499 190 -345 246
rect -289 190 -134 246
rect -78 190 78 246
rect 134 190 289 246
rect 345 190 499 246
rect 555 190 710 246
rect 766 190 921 246
rect 977 190 1132 246
rect 1188 190 1343 246
rect 1399 190 1553 246
rect 1609 190 1764 246
rect 1820 190 1857 246
rect -1857 28 1857 190
rect -1857 -28 -1820 28
rect -1764 -28 -1609 28
rect -1553 -28 -1399 28
rect -1343 -28 -1188 28
rect -1132 -28 -977 28
rect -921 -28 -766 28
rect -710 -28 -555 28
rect -499 -28 -345 28
rect -289 -28 -134 28
rect -78 -28 78 28
rect 134 -28 289 28
rect 345 -28 499 28
rect 555 -28 710 28
rect 766 -28 921 28
rect 977 -28 1132 28
rect 1188 -28 1343 28
rect 1399 -28 1553 28
rect 1609 -28 1764 28
rect 1820 -28 1857 28
rect -1857 -190 1857 -28
rect -1857 -246 -1820 -190
rect -1764 -246 -1609 -190
rect -1553 -246 -1399 -190
rect -1343 -246 -1188 -190
rect -1132 -246 -977 -190
rect -921 -246 -766 -190
rect -710 -246 -555 -190
rect -499 -246 -345 -190
rect -289 -246 -134 -190
rect -78 -246 78 -190
rect 134 -246 289 -190
rect 345 -246 499 -190
rect 555 -246 710 -190
rect 766 -246 921 -190
rect 977 -246 1132 -190
rect 1188 -246 1343 -190
rect 1399 -246 1553 -190
rect 1609 -246 1764 -190
rect 1820 -246 1857 -190
rect -1857 -284 1857 -246
<< properties >>
string GDS_END 1080364
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 1076776
<< end >>
