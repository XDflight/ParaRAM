magic
tech gf180mcuA
timestamp 1666464484
<< properties >>
string GDS_END 256638
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram256x8m8wm1.gds
string GDS_START 256186
<< end >>
