magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< metal1 >>
rect 0 724 1792 844
rect 353 498 399 724
rect 49 60 95 214
rect 801 498 847 724
rect 497 60 543 214
rect 1249 498 1295 724
rect 945 60 991 214
rect 1697 498 1743 724
rect 1393 60 1439 214
rect 0 -60 1792 60
<< obsm1 >>
rect 49 311 95 678
rect 146 392 399 438
rect 49 265 304 311
rect 353 106 399 392
rect 497 311 543 678
rect 594 392 847 438
rect 497 265 752 311
rect 801 106 847 392
rect 945 311 991 678
rect 1042 392 1295 438
rect 945 265 1200 311
rect 1249 106 1295 392
rect 1393 311 1439 678
rect 1490 392 1743 438
rect 1393 265 1648 311
rect 1697 106 1743 392
<< labels >>
rlabel metal1 s 0 724 1792 844 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1697 498 1743 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1249 498 1295 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 801 498 847 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 353 498 399 724 6 VDD
port 1 nsew power bidirectional abutment
rlabel metal1 s 1393 60 1439 214 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 945 60 991 214 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 497 60 543 214 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 49 60 95 214 6 VSS
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -60 1792 60 8 VSS
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1792 784
string LEFclass core SPACER
string LEFsite GF018hv5v_mcu_sc7
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1143332
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/gds/gf180mcu_fd_sc_mcu7t5v0.gds
string GDS_START 1137820
<< end >>
