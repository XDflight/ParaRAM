magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect 4580 2553 5177 2591
rect 3726 2431 5177 2553
rect 2155 2302 5177 2431
rect -532 1217 5177 2302
rect -532 1196 4580 1217
rect -176 1137 4580 1196
rect -176 1096 1540 1137
<< pdiff >>
rect 2814 2062 3097 2290
<< psubdiff >>
rect 3438 2700 3598 2760
rect 3438 2654 3495 2700
rect 3541 2654 3598 2700
rect 3438 2595 3598 2654
rect -352 891 -268 910
rect -352 563 -333 891
rect -287 563 -268 891
rect -352 544 -268 563
rect 4913 -63 4997 -44
rect 4913 -297 4932 -63
rect 4978 -297 4997 -63
rect 4913 -316 4997 -297
<< nsubdiff >>
rect -387 1773 -232 1830
rect -387 1727 -333 1773
rect -287 1727 -232 1773
rect -387 1610 -232 1727
rect -387 1564 -333 1610
rect -287 1564 -232 1610
rect -387 1447 -232 1564
rect -387 1401 -333 1447
rect -287 1401 -232 1447
rect -387 1343 -232 1401
<< psubdiffcont >>
rect 3495 2654 3541 2700
rect -333 563 -287 891
rect 4932 -297 4978 -63
<< nsubdiffcont >>
rect -333 1727 -287 1773
rect -333 1564 -287 1610
rect -333 1401 -287 1447
<< polysilicon >>
rect 2635 2465 2755 2835
rect 3030 2674 3150 2746
rect 4030 2722 4728 2741
rect 4030 2676 4049 2722
rect 4189 2676 4728 2722
rect 4030 2666 4728 2676
rect 4030 2657 4504 2666
rect 3714 2601 3798 2620
rect 2635 2422 2678 2465
rect 2411 2419 2678 2422
rect 2724 2419 2755 2465
rect 3030 2445 3150 2575
rect 3714 2555 3733 2601
rect 3779 2597 3798 2601
rect 3779 2555 4280 2597
rect 3714 2536 4280 2555
rect 3030 2426 3422 2445
rect 3030 2422 3357 2426
rect 2411 2361 2755 2419
rect 3017 2380 3357 2422
rect 3403 2380 3422 2426
rect 3936 2413 4056 2536
rect 4160 2413 4280 2536
rect 4384 2513 4504 2657
rect 4608 2513 4728 2666
rect 3017 2361 3422 2380
rect 3017 2290 3137 2361
rect 3409 1998 3529 2017
rect 3409 1952 3444 1998
rect 3490 1952 3529 1998
rect 79 1166 199 1218
rect 303 1166 423 1218
rect 527 1166 647 1218
rect 751 1166 871 1218
rect 975 1166 1095 1218
rect 1199 1166 1319 1218
rect 79 1147 1521 1166
rect 79 1105 1456 1147
rect 79 968 199 1105
rect 303 968 423 1105
rect 527 968 647 1105
rect 751 968 871 1105
rect 975 968 1095 1105
rect 1199 1101 1456 1105
rect 1502 1101 1521 1147
rect 1199 1082 1521 1101
rect 1199 968 1319 1082
rect 1629 393 1749 1860
rect 2491 1858 3154 1877
rect 3409 1860 3529 1952
rect 2491 1812 3089 1858
rect 3135 1812 3154 1858
rect 2491 1793 3154 1812
rect 2491 1733 2611 1793
rect 2715 1733 2835 1793
rect 2939 1733 3059 1793
rect 3410 1377 3529 1405
rect 2021 1124 2141 1279
rect 1853 1105 2141 1124
rect 1853 1059 1872 1105
rect 2012 1059 2141 1105
rect 1853 1040 2141 1059
rect 2021 480 2141 1040
rect 3409 1028 3529 1377
rect 3410 998 3529 1028
rect 3981 1136 4462 1155
rect 3981 1090 4303 1136
rect 4443 1090 4462 1136
rect 3981 1071 4462 1090
rect 3981 998 4101 1071
rect 4205 998 4325 1071
rect 3410 774 3529 806
rect 2491 484 2611 529
rect 2715 484 2835 529
rect 2939 484 3059 529
rect 3409 511 3529 774
rect 3240 488 3324 507
rect 3240 484 3259 488
rect 2021 461 2214 480
rect 2021 415 2055 461
rect 2195 415 2214 461
rect 2491 442 3259 484
rect 3305 442 3324 488
rect 2491 423 3324 442
rect 3409 492 3588 511
rect 3409 446 3523 492
rect 3569 446 3588 492
rect 3409 427 3588 446
rect 2021 396 2214 415
rect 1597 374 1775 393
rect 1597 328 1616 374
rect 1756 328 1775 374
rect 1597 309 1775 328
rect 4429 216 4549 360
rect 4653 216 4773 360
rect 4429 197 4773 216
rect 4429 151 4525 197
rect 4665 151 4773 197
rect 4429 132 4773 151
<< polycontact >>
rect 4049 2676 4189 2722
rect 2678 2419 2724 2465
rect 3733 2555 3779 2601
rect 3357 2380 3403 2426
rect 3444 1952 3490 1998
rect 1456 1101 1502 1147
rect 3089 1812 3135 1858
rect 1872 1059 2012 1105
rect 4303 1090 4443 1136
rect 2055 415 2195 461
rect 3259 442 3305 488
rect 3523 446 3569 492
rect 1616 328 1756 374
rect 4525 151 4665 197
<< metal1 >>
rect 2784 2853 2941 3324
rect 2784 2778 3519 2853
rect -367 1773 -252 1810
rect -367 1727 -333 1773
rect -287 1727 -252 1773
rect -367 1610 -252 1727
rect 194 1665 310 2191
rect 642 1665 758 2191
rect 1124 1665 1170 2239
rect 2170 2005 2216 2713
rect 2560 1923 2606 2753
rect 2784 2553 3001 2778
rect 3447 2751 3519 2778
rect 3709 2790 3801 2830
rect 3447 2700 3589 2751
rect 3131 2476 3247 2699
rect 3447 2654 3495 2700
rect 3541 2654 3589 2700
rect 3447 2604 3589 2654
rect 3709 2738 3729 2790
rect 3781 2738 3801 2790
rect 3709 2604 3801 2738
rect 4038 2722 4200 2733
rect 4038 2676 4049 2722
rect 4189 2676 4200 2722
rect 4038 2665 4200 2676
rect 3709 2552 3729 2604
rect 3781 2552 3801 2604
rect 3709 2511 3801 2552
rect 3861 2563 4803 2609
rect 2667 2465 3247 2476
rect 2667 2419 2678 2465
rect 2724 2419 3247 2465
rect 2667 2402 3247 2419
rect 3131 2152 3247 2402
rect 3324 2426 3580 2445
rect 3861 2435 3907 2563
rect 3324 2380 3357 2426
rect 3403 2415 3580 2426
rect 3324 2363 3363 2380
rect 3415 2363 3580 2415
rect 4309 2413 4355 2563
rect 4757 2435 4803 2563
rect 3324 2290 3580 2363
rect 3263 2023 3602 2064
rect 3263 2004 3300 2023
rect 3098 1971 3300 2004
rect 3352 1998 3512 2023
rect 3352 1971 3444 1998
rect 3098 1952 3444 1971
rect 3490 1971 3512 1998
rect 3564 1971 3602 2023
rect 3490 1952 3602 1971
rect 3098 1929 3602 1952
rect 2382 1804 2946 1923
rect 3098 1869 3170 1929
rect -367 1564 -333 1610
rect -287 1564 -252 1610
rect -367 1447 -252 1564
rect -367 1401 -333 1447
rect -287 1401 -252 1447
rect -367 1364 -252 1401
rect 4 1166 50 1445
rect 452 1166 498 1445
rect 900 1166 946 1445
rect 1348 1166 1394 1445
rect 4 1046 1394 1166
rect 1468 1158 1648 1166
rect 1445 1154 1648 1158
rect 1445 1147 1480 1154
rect 1445 1101 1456 1147
rect 1636 1102 1648 1154
rect 1502 1101 1648 1102
rect 1445 1090 1648 1101
rect 1778 1116 1824 1315
rect 1778 1105 2023 1116
rect -344 891 -276 902
rect -344 563 -333 891
rect -287 563 -276 891
rect 4 779 50 1046
rect -344 552 -276 563
rect 194 348 310 901
rect 452 779 498 1046
rect 642 348 758 901
rect 900 779 946 1046
rect 1090 348 1206 901
rect 1348 779 1394 1046
rect 1778 1059 1872 1105
rect 2012 1059 2023 1105
rect 1778 1048 2023 1059
rect 1778 798 1824 1048
rect 2170 798 2216 1315
rect 2382 544 2498 1804
rect 2160 472 2206 476
rect 2044 461 2206 472
rect 2044 415 2055 461
rect 2195 415 2206 461
rect 2044 404 2206 415
rect 1600 376 1780 388
rect 1600 324 1612 376
rect 1768 324 1780 376
rect 1600 312 1780 324
rect 2160 237 2206 404
rect 2606 472 2722 1722
rect 2830 544 2946 1804
rect 3078 1858 3170 1869
rect 3078 1812 3089 1858
rect 3135 1812 3170 1858
rect 3078 1801 3170 1812
rect 3054 472 3170 1724
rect 3334 863 3380 1803
rect 4085 1194 4131 1424
rect 3951 1182 4131 1194
rect 3951 1130 3963 1182
rect 4119 1130 4131 1182
rect 3951 1118 4131 1130
rect 3282 807 3380 863
rect 4085 957 4131 1118
rect 4280 1139 4460 1151
rect 4280 1087 4292 1139
rect 4448 1087 4460 1139
rect 4280 1075 4460 1087
rect 4085 862 4161 957
rect 3282 499 3354 807
rect 2606 353 3170 472
rect 3248 488 3354 499
rect 3248 442 3259 488
rect 3305 442 3354 488
rect 3248 432 3354 442
rect 3432 493 3771 534
rect 3432 441 3469 493
rect 3521 492 3681 493
rect 3521 446 3523 492
rect 3569 446 3681 492
rect 3521 441 3681 446
rect 3733 441 3771 493
rect 3248 431 3316 432
rect 3432 400 3771 441
rect 3906 330 3952 463
rect 4354 330 4400 485
rect 4802 330 4848 463
rect 3906 284 4848 330
rect 2160 197 3783 237
rect 4514 197 4676 208
rect 2160 191 4525 197
rect 3702 151 4525 191
rect 4665 151 4676 197
rect 4514 140 4676 151
rect 4921 -63 4989 -52
rect 4921 -297 4932 -63
rect 4978 -297 4989 -63
rect 4921 -308 4989 -297
<< via1 >>
rect 3729 2738 3781 2790
rect 3729 2601 3781 2604
rect 3729 2555 3733 2601
rect 3733 2555 3779 2601
rect 3779 2555 3781 2601
rect 3729 2552 3781 2555
rect 3363 2380 3403 2415
rect 3403 2380 3415 2415
rect 3363 2363 3415 2380
rect 3300 1971 3352 2023
rect 3512 1971 3564 2023
rect 1480 1147 1636 1154
rect 1480 1102 1502 1147
rect 1502 1102 1636 1147
rect 1612 374 1768 376
rect 1612 328 1616 374
rect 1616 328 1756 374
rect 1756 328 1768 374
rect 1612 324 1768 328
rect 3963 1130 4119 1182
rect 4292 1136 4448 1139
rect 4292 1090 4303 1136
rect 4303 1090 4443 1136
rect 4443 1090 4448 1136
rect 4292 1087 4448 1090
rect 3469 441 3521 493
rect 3681 441 3733 493
<< metal2 >>
rect 3709 2790 3801 2830
rect 3709 2751 3729 2790
rect 3708 2738 3729 2751
rect 3781 2751 3801 2790
rect 3781 2738 3802 2751
rect 3708 2604 3802 2738
rect 3708 2552 3729 2604
rect 3781 2552 3802 2604
rect 3076 2415 3452 2438
rect 3076 2363 3363 2415
rect 3415 2363 3452 2415
rect 3076 2341 3452 2363
rect 1468 1165 1648 1166
rect 1468 1155 1671 1165
rect 1468 1154 1501 1155
rect 1468 1102 1480 1154
rect 1468 1099 1501 1102
rect 1661 1099 1671 1155
rect 3076 1103 3170 2341
rect 3263 2023 3602 2064
rect 3263 1971 3300 2023
rect 3352 1971 3512 2023
rect 3564 1971 3602 2023
rect 3263 1930 3602 1971
rect 1468 1090 1671 1099
rect 1491 1089 1671 1090
rect 3344 534 3433 1930
rect 3708 1060 3802 2552
rect 3951 1184 4131 1194
rect 3951 1128 3961 1184
rect 4121 1128 4131 1184
rect 4324 1151 4418 2751
rect 3951 1118 4131 1128
rect 4280 1139 4460 1151
rect 4280 1087 4292 1139
rect 4448 1087 4460 1139
rect 4280 1075 4460 1087
rect 3344 493 3771 534
rect 3344 441 3469 493
rect 3521 441 3681 493
rect 3733 441 3771 493
rect 3344 400 3771 441
rect 1600 376 1780 388
rect 1600 324 1612 376
rect 1768 324 1780 376
rect 1600 312 1780 324
<< via2 >>
rect 1501 1154 1661 1155
rect 1501 1102 1636 1154
rect 1636 1102 1661 1154
rect 1501 1099 1661 1102
rect 3961 1182 4121 1184
rect 3961 1130 3963 1182
rect 3963 1130 4119 1182
rect 4119 1130 4121 1182
rect 3961 1128 4121 1130
<< metal3 >>
rect 2113 2655 4296 2748
rect -356 1502 5006 2312
rect 1491 1184 4131 1203
rect 1491 1155 3961 1184
rect 1491 1099 1501 1155
rect 1661 1128 3961 1155
rect 4121 1128 4131 1184
rect 1661 1106 4131 1128
rect 1661 1099 1671 1106
rect 1491 1089 1671 1099
rect -356 169 5028 957
rect -357 -359 5028 169
use M1_NACTIVE4310591302038_512x8m81  M1_NACTIVE4310591302038_512x8m81_0
timestamp 1666464484
transform 1 0 4955 0 1 1951
box -42 -418 42 418
use M1_NACTIVE4310591302041_512x8m81  M1_NACTIVE4310591302041_512x8m81_0
timestamp 1666464484
transform 1 0 478 0 1 2177
box -700 -42 700 42
use M1_NWELL_01_R270_512x8m81  M1_NWELL_01_R270_512x8m81_0
timestamp 1666464484
transform 0 1 -310 -1 0 1587
box 0 0 1 1
use M1_PACTIVE4310591302034_512x8m81  M1_PACTIVE4310591302034_512x8m81_0
timestamp 1666464484
transform 1 0 -310 0 1 727
box 0 0 1 1
use M1_PACTIVE4310591302039_512x8m81  M1_PACTIVE4310591302039_512x8m81_0
timestamp 1666464484
transform 1 0 4955 0 1 -180
box 0 0 1 1
use M1_PACTIVE4310591302040_512x8m81  M1_PACTIVE4310591302040_512x8m81_0
timestamp 1666464484
transform 1 0 683 0 1 338
box -747 -42 747 42
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_0
timestamp 1666464484
transform 0 -1 1479 1 0 1124
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_1
timestamp 1666464484
transform 1 0 3546 0 1 469
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_2
timestamp 1666464484
transform 1 0 2701 0 1 2442
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_3
timestamp 1666464484
transform 1 0 3380 0 1 2403
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_4
timestamp 1666464484
transform 1 0 3112 0 1 1835
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_5
timestamp 1666464484
transform 1 0 3467 0 1 1975
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_6
timestamp 1666464484
transform 1 0 3756 0 1 2578
box 0 0 1 1
use M1_POLY24310591302031_512x8m81  M1_POLY24310591302031_512x8m81_7
timestamp 1666464484
transform 1 0 3282 0 1 465
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_0
timestamp 1666464484
transform -1 0 2125 0 -1 438
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_1
timestamp 1666464484
transform -1 0 1942 0 -1 1082
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_2
timestamp 1666464484
transform 1 0 4119 0 -1 2699
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_3
timestamp 1666464484
transform 1 0 4595 0 1 174
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_4
timestamp 1666464484
transform 1 0 1686 0 1 351
box 0 0 1 1
use M1_POLY24310591302033_512x8m81  M1_POLY24310591302033_512x8m81_5
timestamp 1666464484
transform 1 0 4373 0 1 1113
box 0 0 1 1
use M1_PSUB_02_512x8m81  M1_PSUB_02_512x8m81_0
timestamp 1666464484
transform 1 0 3518 0 1 2677
box 0 0 1 1
use M2_M1$$168351788_R90_512x8m81  M2_M1$$168351788_R90_512x8m81_0
timestamp 1666464484
transform 0 -1 3601 1 0 467
box 0 0 1 1
use M2_M1$$168351788_R90_512x8m81  M2_M1$$168351788_R90_512x8m81_1
timestamp 1666464484
transform 0 -1 3432 1 0 1997
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_0
timestamp 1666464484
transform 1 0 1690 0 1 350
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_1
timestamp 1666464484
transform 1 0 1558 0 1 1128
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_2
timestamp 1666464484
transform 1 0 4041 0 1 1156
box 0 0 1 1
use M2_M1431059130200_512x8m81  M2_M1431059130200_512x8m81_3
timestamp 1666464484
transform 1 0 4370 0 1 1113
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_0
timestamp 1666464484
transform 1 0 4041 0 1 1156
box 0 0 1 1
use M3_M2431059130207_512x8m81  M3_M2431059130207_512x8m81_1
timestamp 1666464484
transform 1 0 1581 0 1 1127
box 0 0 1 1
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_0
timestamp 1666464484
transform -1 0 3529 0 1 807
box -88 -44 208 236
use nmos_5p0431059130208_512x8m81  nmos_5p0431059130208_512x8m81_1
timestamp 1666464484
transform 1 0 2635 0 -1 2761
box -88 -44 208 236
use nmos_5p04310591302033_512x8m81  nmos_5p04310591302033_512x8m81_0
timestamp 1666464484
transform 1 0 3030 0 -1 2673
box -88 -44 208 164
use nmos_5p04310591302044_512x8m81  nmos_5p04310591302044_512x8m81_0
timestamp 1666464484
transform -1 0 2141 0 1 540
box -88 -44 208 484
use nmos_5p04310591302045_512x8m81  nmos_5p04310591302045_512x8m81_0
timestamp 1666464484
transform 1 0 4429 0 -1 957
box -88 -44 432 612
use nmos_5p04310591302045_512x8m81  nmos_5p04310591302045_512x8m81_1
timestamp 1666464484
transform 1 0 3981 0 -1 957
box -88 -44 432 612
use nmos_5p04310591302046_512x8m81  nmos_5p04310591302046_512x8m81_0
timestamp 1666464484
transform -1 0 1319 0 -1 957
box -88 -44 1328 468
use nmos_5p04310591302050_512x8m81  nmos_5p04310591302050_512x8m81_0
timestamp 1666464484
transform -1 0 3059 0 1 544
box -88 -44 656 498
use nmos_5p04310591302052_512x8m81  nmos_5p04310591302052_512x8m81_0
timestamp 1666464484
transform -1 0 1749 0 1 544
box -88 -44 208 364
use pmos_1p2$$171625516_512x8m81  pmos_1p2$$171625516_512x8m81_0
timestamp 1666464484
transform 1 0 2442 0 -1 2290
box -286 -142 568 348
use pmos_5p04310591302013_512x8m81  pmos_5p04310591302013_512x8m81_0
timestamp 1666464484
transform -1 0 3059 0 1 1279
box -208 -120 776 574
use pmos_5p04310591302014_512x8m81  pmos_5p04310591302014_512x8m81_0
timestamp 1666464484
transform -1 0 3529 0 1 1406
box -208 -120 328 574
use pmos_5p04310591302038_512x8m81  pmos_5p04310591302038_512x8m81_0
timestamp 1666464484
transform 1 0 3017 0 -1 2290
box -208 -120 328 360
use pmos_5p04310591302047_512x8m81  pmos_5p04310591302047_512x8m81_0
timestamp 1666464484
transform -1 0 1749 0 1 1279
box -208 -120 328 920
use pmos_5p04310591302048_512x8m81  pmos_5p04310591302048_512x8m81_0
timestamp 1666464484
transform -1 0 2141 0 1 1235
box -208 -120 328 1020
use pmos_5p04310591302049_512x8m81  pmos_5p04310591302049_512x8m81_0
timestamp 1666464484
transform -1 0 1319 0 1 1238
box -208 -120 1448 876
use pmos_5p04310591302051_512x8m81  pmos_5p04310591302051_512x8m81_0
timestamp 1666464484
transform 1 0 3936 0 1 1337
box -208 -120 552 1254
use pmos_5p04310591302051_512x8m81  pmos_5p04310591302051_512x8m81_1
timestamp 1666464484
transform 1 0 4384 0 1 1337
box -208 -120 552 1254
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_0
timestamp 1666464484
transform -1 0 3169 0 1 1086
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_1
timestamp 1666464484
transform -1 0 2710 0 1 1086
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_2
timestamp 1666464484
transform 0 -1 4226 1 0 2655
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_3
timestamp 1666464484
transform 0 -1 2478 1 0 2655
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_4
timestamp 1666464484
transform 1 0 4909 0 1 -340
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_5
timestamp 1666464484
transform 1 0 206 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_6
timestamp 1666464484
transform 1 0 652 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_7
timestamp 1666464484
transform 1 0 1100 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_8
timestamp 1666464484
transform 1 0 652 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_9
timestamp 1666464484
transform 1 0 206 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_10
timestamp 1666464484
transform 1 0 4510 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_11
timestamp 1666464484
transform 1 0 4510 0 1 2004
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_12
timestamp 1666464484
transform 1 0 4555 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_13
timestamp 1666464484
transform 1 0 3525 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_14
timestamp 1666464484
transform 1 0 3547 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_15
timestamp 1666464484
transform 1 0 1102 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_16
timestamp 1666464484
transform 1 0 2761 0 1 2004
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_17
timestamp 1666464484
transform 1 0 2312 0 1 2004
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_18
timestamp 1666464484
transform 1 0 -356 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_19
timestamp 1666464484
transform 1 0 -356 0 1 630
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_20
timestamp 1666464484
transform 1 0 4909 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_21
timestamp 1666464484
transform 1 0 4909 0 1 2004
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_22
timestamp 1666464484
transform 1 0 1531 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_23
timestamp 1666464484
transform 1 0 1923 0 1 1503
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_24
timestamp 1666464484
transform 1 0 1531 0 1 537
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_25
timestamp 1666464484
transform 1 0 1923 0 1 537
box 0 -1 93 308
use via1_2_x2_512x8m81  via1_2_x2_512x8m81_26
timestamp 1666464484
transform 1 0 2919 0 1 2004
box 0 -1 93 308
use via1_R270_512x8m81  via1_R270_512x8m81_0
timestamp 1666464484
transform 0 1 3325 -1 0 2437
box 0 0 1 1
use via1_x2_512x8m81  via1_x2_512x8m81_0
timestamp 1666464484
transform -1 0 3801 0 1 2512
box 0 0 1 1
<< labels >>
rlabel metal3 s -214 644 -214 644 4 vss
port 1 nsew
rlabel metal3 s -255 2131 -255 2131 4 vdd
port 2 nsew
rlabel metal2 s 3762 2693 3762 2693 4 qp
port 3 nsew
rlabel metal2 s 4401 2693 4401 2693 4 qn
port 4 nsew
rlabel metal1 s 3628 469 3628 469 4 se
port 5 nsew
rlabel metal1 s 467 1145 467 1145 4 q
port 6 nsew
rlabel metal1 s 3511 2689 3511 2689 4 vss
port 1 nsew
rlabel metal1 s 1613 361 1613 361 4 GWE
port 7 nsew
<< properties >>
string GDS_END 421544
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 410570
string path 21.660 12.815 21.660 12.970 
<< end >>
