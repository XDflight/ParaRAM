magic
tech gf180mcuA
magscale 1 10
timestamp 1666464484
<< polysilicon >>
rect -31 567 89 640
rect 193 567 313 640
rect 417 567 537 640
rect 641 567 761 640
rect 865 567 985 640
rect 1089 567 1209 640
rect 1313 567 1433 640
rect 1537 567 1657 640
rect -31 -74 89 -1
rect 193 -74 313 -1
rect 417 -74 537 -1
rect 641 -74 761 -1
rect 865 -74 985 -1
rect 1089 -74 1209 -1
rect 1313 -74 1433 -1
rect 1537 -74 1657 -1
use nmos_5p04310591302017_512x8m81  nmos_5p04310591302017_512x8m81_0
timestamp 1666464484
transform 1 0 -31 0 1 0
box -88 -44 1776 612
<< properties >>
string GDS_END 258286
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram512x8m8wm1.gds
string GDS_START 257140
<< end >>
