magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< mvnmos >>
rect 0 0 200 120
<< mvndiff >>
rect -88 83 0 120
rect -88 37 -75 83
rect -29 37 0 83
rect -88 0 0 37
rect 200 83 288 120
rect 200 37 229 83
rect 275 37 288 83
rect 200 0 288 37
<< mvndiffc >>
rect -75 37 -29 83
rect 229 37 275 83
<< polysilicon >>
rect 0 120 200 164
rect 0 -44 200 0
<< metal1 >>
rect -75 83 -29 120
rect -75 0 -29 37
rect 229 83 275 120
rect 229 0 275 37
<< labels >>
flabel metal1 s -52 60 -52 60 0 FreeSans 200 0 0 0 S
flabel metal1 s 252 60 252 60 0 FreeSans 200 0 0 0 D
<< properties >>
string GDS_END 922972
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_ip_sram/gds/gf180mcu_fd_ip_sram__sram64x8m8wm1.gds
string GDS_START 921948
<< end >>
