magic
tech gf180mcuB
magscale 1 10
timestamp 1666464484
<< nwell >>
rect -86 453 3446 1094
<< pwell >>
rect -86 -86 3446 453
<< mvnmos >>
rect 124 156 244 296
rect 348 156 468 296
rect 572 156 692 296
rect 796 156 916 296
rect 1012 156 1132 296
rect 1236 156 1356 296
rect 1604 157 1724 297
rect 1828 157 1948 297
rect 2284 157 2404 297
rect 2508 157 2628 297
rect 2732 157 2852 297
rect 3100 123 3220 323
<< mvpmos >>
rect 210 576 310 852
rect 358 576 458 852
rect 582 576 682 852
rect 884 576 984 852
rect 1032 576 1132 852
rect 1236 576 1336 852
rect 1604 573 1704 849
rect 1808 573 1908 849
rect 2320 573 2420 849
rect 2524 573 2624 849
rect 2672 573 2772 849
rect 3110 573 3210 939
<< mvndiff >>
rect 36 216 124 296
rect 36 170 49 216
rect 95 170 124 216
rect 36 156 124 170
rect 244 216 348 296
rect 244 170 273 216
rect 319 170 348 216
rect 244 156 348 170
rect 468 216 572 296
rect 468 170 497 216
rect 543 170 572 216
rect 468 156 572 170
rect 692 216 796 296
rect 692 170 721 216
rect 767 170 796 216
rect 692 156 796 170
rect 916 156 1012 296
rect 1132 216 1236 296
rect 1132 170 1161 216
rect 1207 170 1236 216
rect 1132 156 1236 170
rect 1356 216 1444 296
rect 1356 170 1385 216
rect 1431 170 1444 216
rect 1356 156 1444 170
rect 1516 216 1604 297
rect 1516 170 1529 216
rect 1575 170 1604 216
rect 1516 157 1604 170
rect 1724 216 1828 297
rect 1724 170 1753 216
rect 1799 170 1828 216
rect 1724 157 1828 170
rect 1948 216 2036 297
rect 1948 170 1977 216
rect 2023 170 2036 216
rect 1948 157 2036 170
rect 3012 310 3100 323
rect 2196 216 2284 297
rect 2196 170 2209 216
rect 2255 170 2284 216
rect 2196 157 2284 170
rect 2404 216 2508 297
rect 2404 170 2433 216
rect 2479 170 2508 216
rect 2404 157 2508 170
rect 2628 216 2732 297
rect 2628 170 2657 216
rect 2703 170 2732 216
rect 2628 157 2732 170
rect 2852 216 2940 297
rect 2852 170 2881 216
rect 2927 170 2940 216
rect 2852 157 2940 170
rect 3012 170 3025 310
rect 3071 170 3100 310
rect 3012 123 3100 170
rect 3220 310 3308 323
rect 3220 170 3249 310
rect 3295 170 3308 310
rect 3220 123 3308 170
<< mvpdiff >>
rect 122 829 210 852
rect 122 689 135 829
rect 181 689 210 829
rect 122 576 210 689
rect 310 576 358 852
rect 458 576 582 852
rect 682 829 884 852
rect 682 689 711 829
rect 757 689 884 829
rect 682 576 884 689
rect 984 576 1032 852
rect 1132 829 1236 852
rect 1132 689 1161 829
rect 1207 689 1236 829
rect 1132 576 1236 689
rect 1336 769 1424 852
rect 1336 629 1365 769
rect 1411 629 1424 769
rect 1336 576 1424 629
rect 1516 769 1604 849
rect 1516 629 1529 769
rect 1575 629 1604 769
rect 1516 573 1604 629
rect 1704 829 1808 849
rect 1704 689 1733 829
rect 1779 689 1808 829
rect 1704 573 1808 689
rect 1908 829 1996 849
rect 1908 689 1937 829
rect 1983 689 1996 829
rect 1908 573 1996 689
rect 2232 769 2320 849
rect 2232 629 2245 769
rect 2291 629 2320 769
rect 2232 573 2320 629
rect 2420 829 2524 849
rect 2420 689 2449 829
rect 2495 689 2524 829
rect 2420 573 2524 689
rect 2624 573 2672 849
rect 2772 829 2860 849
rect 2772 689 2801 829
rect 2847 689 2860 829
rect 2772 573 2860 689
rect 3022 829 3110 939
rect 3022 689 3035 829
rect 3081 689 3110 829
rect 3022 573 3110 689
rect 3210 829 3298 939
rect 3210 689 3239 829
rect 3285 689 3298 829
rect 3210 573 3298 689
<< mvndiffc >>
rect 49 170 95 216
rect 273 170 319 216
rect 497 170 543 216
rect 721 170 767 216
rect 1161 170 1207 216
rect 1385 170 1431 216
rect 1529 170 1575 216
rect 1753 170 1799 216
rect 1977 170 2023 216
rect 2209 170 2255 216
rect 2433 170 2479 216
rect 2657 170 2703 216
rect 2881 170 2927 216
rect 3025 170 3071 310
rect 3249 170 3295 310
<< mvpdiffc >>
rect 135 689 181 829
rect 711 689 757 829
rect 1161 689 1207 829
rect 1365 629 1411 769
rect 1529 629 1575 769
rect 1733 689 1779 829
rect 1937 689 1983 829
rect 2245 629 2291 769
rect 2449 689 2495 829
rect 2801 689 2847 829
rect 3035 689 3081 829
rect 3239 689 3285 829
<< polysilicon >>
rect 1032 944 1908 984
rect 210 852 310 896
rect 358 852 458 896
rect 582 852 682 896
rect 884 852 984 896
rect 1032 852 1132 944
rect 1236 852 1336 896
rect 1604 849 1704 893
rect 1808 849 1908 944
rect 3110 939 3210 983
rect 2320 849 2420 893
rect 2524 849 2624 893
rect 2672 849 2772 893
rect 210 532 310 576
rect 210 455 250 532
rect 124 442 250 455
rect 124 396 137 442
rect 183 433 250 442
rect 358 442 458 576
rect 582 516 682 576
rect 884 540 984 576
rect 582 476 836 516
rect 884 494 897 540
rect 943 494 984 540
rect 884 481 984 494
rect 183 396 244 433
rect 124 296 244 396
rect 358 396 371 442
rect 417 396 458 442
rect 358 340 458 396
rect 572 415 748 428
rect 572 369 689 415
rect 735 369 748 415
rect 572 356 748 369
rect 348 296 468 340
rect 572 296 692 356
rect 796 340 836 476
rect 1032 340 1132 576
rect 796 296 916 340
rect 1012 296 1132 340
rect 1236 340 1336 576
rect 1604 442 1704 573
rect 1604 396 1621 442
rect 1667 396 1704 442
rect 1604 341 1704 396
rect 1808 442 1908 573
rect 2320 529 2420 573
rect 2320 455 2404 529
rect 1808 396 1821 442
rect 1867 396 1908 442
rect 1808 383 1908 396
rect 2064 442 2136 455
rect 2064 396 2077 442
rect 2123 396 2136 442
rect 2064 383 2136 396
rect 1828 341 1908 383
rect 1236 296 1356 340
rect 1604 297 1724 341
rect 1828 297 1948 341
rect 124 112 244 156
rect 348 112 468 156
rect 572 112 692 156
rect 796 112 916 156
rect 1012 112 1132 156
rect 876 64 916 112
rect 1236 64 1356 156
rect 1604 113 1724 157
rect 1828 113 1948 157
rect 2096 64 2136 383
rect 2284 442 2404 455
rect 2284 396 2297 442
rect 2343 396 2404 442
rect 2284 297 2404 396
rect 2524 442 2624 573
rect 2672 529 2772 573
rect 2524 396 2537 442
rect 2583 396 2624 442
rect 2524 341 2624 396
rect 2732 341 2772 529
rect 3110 455 3210 573
rect 3078 442 3210 455
rect 3078 396 3091 442
rect 3137 396 3210 442
rect 3078 383 3210 396
rect 3100 367 3210 383
rect 2508 297 2628 341
rect 2732 297 2852 341
rect 3100 323 3220 367
rect 876 24 2136 64
rect 2284 65 2404 157
rect 2508 113 2628 157
rect 2732 65 2852 157
rect 3100 79 3220 123
rect 2284 25 2852 65
<< polycontact >>
rect 137 396 183 442
rect 897 494 943 540
rect 371 396 417 442
rect 689 369 735 415
rect 1621 396 1667 442
rect 1821 396 1867 442
rect 2077 396 2123 442
rect 2297 396 2343 442
rect 2537 396 2583 442
rect 3091 396 3137 442
<< metal1 >>
rect 0 918 3360 1098
rect 135 829 181 918
rect 135 678 181 689
rect 711 829 757 840
rect 711 632 757 689
rect 1161 829 1207 918
rect 1161 678 1207 689
rect 1253 826 1667 872
rect 1253 632 1299 826
rect 597 586 1299 632
rect 1365 769 1431 780
rect 1411 629 1431 769
rect 30 453 82 542
rect 30 442 183 453
rect 30 396 137 442
rect 30 354 183 396
rect 242 442 418 453
rect 242 396 371 442
rect 417 396 418 442
rect 242 354 418 396
rect 49 262 543 308
rect 49 216 95 262
rect 497 216 543 262
rect 49 159 95 170
rect 262 170 273 216
rect 319 170 330 216
rect 262 90 330 170
rect 597 216 643 586
rect 1365 540 1431 629
rect 689 494 897 540
rect 943 494 1431 540
rect 689 415 735 494
rect 689 358 735 369
rect 1161 216 1207 227
rect 597 170 721 216
rect 767 170 778 216
rect 497 159 543 170
rect 1161 90 1207 170
rect 1385 216 1431 494
rect 1385 159 1431 170
rect 1529 769 1575 780
rect 1529 339 1575 629
rect 1621 442 1667 826
rect 1733 829 1779 918
rect 1733 678 1779 689
rect 1937 829 2403 872
rect 1983 826 2403 829
rect 1983 689 2023 826
rect 1621 385 1667 396
rect 1713 396 1821 442
rect 1867 396 1878 442
rect 1713 339 1759 396
rect 1529 293 1759 339
rect 1529 216 1575 293
rect 1529 159 1575 170
rect 1753 216 1799 227
rect 1753 90 1799 170
rect 1937 216 2023 689
rect 2245 769 2291 780
rect 1937 170 1977 216
rect 2077 629 2245 634
rect 2077 588 2291 629
rect 2357 632 2403 826
rect 2449 829 2495 918
rect 2449 678 2495 689
rect 2801 829 2847 840
rect 2077 442 2123 588
rect 2357 586 2583 632
rect 2077 216 2123 396
rect 2270 442 2343 542
rect 2270 396 2297 442
rect 2270 354 2343 396
rect 2537 442 2583 586
rect 2537 385 2583 396
rect 2801 442 2847 689
rect 3035 829 3081 918
rect 3239 829 3295 840
rect 3035 678 3081 689
rect 3166 689 3239 766
rect 3285 689 3295 829
rect 3166 678 3295 689
rect 2801 396 3091 442
rect 3137 396 3148 442
rect 2801 304 2847 396
rect 2657 258 2847 304
rect 3025 310 3071 321
rect 3249 318 3295 678
rect 2433 216 2479 227
rect 2077 170 2209 216
rect 2255 170 2266 216
rect 1937 159 2023 170
rect 2433 90 2479 170
rect 2657 216 2703 258
rect 2657 159 2703 170
rect 2881 216 2927 227
rect 2881 90 2927 170
rect 3166 310 3295 318
rect 3166 242 3249 310
rect 3025 90 3071 170
rect 3249 159 3295 170
rect 0 -90 3360 90
<< labels >>
flabel metal1 s 2270 354 2343 542 0 FreeSans 200 0 0 0 CLKN
port 1 nsew clock input
flabel metal1 s 242 354 418 453 0 FreeSans 200 0 0 0 E
port 2 nsew default input
flabel metal1 s 3239 766 3295 840 0 FreeSans 200 0 0 0 Q
port 4 nsew default output
flabel metal1 s 30 453 82 542 0 FreeSans 200 0 0 0 TE
port 3 nsew default input
flabel metal1 s 0 918 3360 1098 0 FreeSans 200 0 0 0 VDD
port 5 nsew power bidirectional abutment
flabel metal1 s 3025 227 3071 321 0 FreeSans 200 0 0 0 VSS
port 8 nsew ground bidirectional abutment
flabel pwell 0 400 0 400 3 FreeSans 600 0 0 0 & Vendor GLOBALFOUNDRIES
flabel pwell 0 300 0 300 3 FreeSans 600 0 0 0 & Product GF018hv5v_green_sc9
flabel pwell 0 200 0 200 3 FreeSans 600 0 0 0 & Version 2015q2v2
flabel pwell 0 100 0 100 3 FreeSans 600 0 0 0 & Metric 1.00
rlabel metal1 s 30 354 183 453 1 TE
port 3 nsew default input
rlabel metal1 s 3166 678 3295 766 1 Q
port 4 nsew default output
rlabel metal1 s 3249 318 3295 678 1 Q
port 4 nsew default output
rlabel metal1 s 3166 242 3295 318 1 Q
port 4 nsew default output
rlabel metal1 s 3249 159 3295 242 1 Q
port 4 nsew default output
rlabel metal1 s 3035 678 3081 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 2449 678 2495 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1733 678 1779 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 1161 678 1207 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 135 678 181 918 1 VDD
port 5 nsew power bidirectional abutment
rlabel metal1 s 3025 216 3071 227 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2881 216 2927 227 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2433 216 2479 227 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1753 216 1799 227 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1161 216 1207 227 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 3025 90 3071 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2881 90 2927 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 2433 90 2479 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1753 90 1799 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 1161 90 1207 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 262 90 330 216 1 VSS
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 -90 3360 90 1 VSS
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 3360 1008
string GDS_END 811424
string GDS_FILE $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu9t5v0/gds/gf180mcu_fd_sc_mcu9t5v0.gds
string GDS_START 803628
string LEFclass core
string LEFsite GF018hv5v_green_sc9
string LEFsymmetry X Y
<< end >>
